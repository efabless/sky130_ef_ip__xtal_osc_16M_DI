VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_16M_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_16M_DI ;
  ORIGIN -70.855 0.000 ;
  SIZE 454.445 BY 211.800 ;
  PIN dout
    ANTENNADIFFAREA 0.435000 ;
    PORT
      LAYER met2 ;
        RECT 213.640 -3.280 213.920 60.465 ;
    END
  END dout
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER met2 ;
        RECT 519.780 134.970 520.420 218.525 ;
    END
  END in
  PIN ena
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER met2 ;
        RECT 208.390 -3.280 208.670 61.955 ;
    END
  END ena
  PIN stdby
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER met2 ;
        RECT 221.075 -3.280 221.355 62.785 ;
    END
  END stdby
  PIN out
    PORT
      LAYER met2 ;
        RECT 74.780 134.970 75.420 218.525 ;
    END
  END out
  PIN vssd1
    ANTENNADIFFAREA 21.305099 ;
    PORT
      LAYER met4 ;
        RECT 187.275 0.000 188.875 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 192.605 0.000 194.205 211.800 ;
    END
  END vssd1
  PIN vdda1
    ANTENNADIFFAREA 98.890800 ;
    PORT
      LAYER met4 ;
        RECT 226.550 0.000 228.150 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 222.405 0.000 224.005 211.800 ;
    END
  END vdda1
  PIN vccd1
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER met4 ;
        RECT 216.610 0.000 218.210 211.800 ;
    END
  END vccd1
  PIN vssa1
    ANTENNADIFFAREA 81.684601 ;
    PORT
      LAYER met4 ;
        RECT 206.090 0.000 207.690 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.565 0.000 203.165 211.800 ;
    END
  END vssa1
  OBS
      LAYER li1 ;
        RECT 201.420 62.550 229.015 116.595 ;
      LAYER met1 ;
        RECT 185.745 60.240 229.045 117.060 ;
      LAYER met2 ;
        RECT 75.700 134.690 519.500 135.970 ;
        RECT 75.420 63.065 519.780 134.690 ;
        RECT 75.420 62.235 220.795 63.065 ;
        RECT 75.420 0.000 208.110 62.235 ;
        RECT 208.950 60.745 220.795 62.235 ;
        RECT 208.950 0.000 213.360 60.745 ;
        RECT 214.200 0.000 220.795 60.745 ;
        RECT 221.635 0.000 519.780 63.065 ;
      LAYER met3 ;
        RECT 186.875 62.420 229.275 117.060 ;
  END
END sky130_ef_ip__xtal_osc_16M_DI
END LIBRARY

