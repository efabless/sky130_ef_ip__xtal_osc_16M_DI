VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_16M_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_16M_DI ;
  ORIGIN -70.855 0.000 ;
  SIZE 454.445 BY 211.800 ;
  PIN dout
    ANTENNADIFFAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 214.180 64.640 214.350 65.180 ;
        RECT 216.110 63.650 216.280 64.690 ;
      LAYER mcon ;
        RECT 214.180 64.825 214.350 64.995 ;
        RECT 216.110 64.265 216.280 64.435 ;
        RECT 216.110 63.905 216.280 64.075 ;
      LAYER met1 ;
        RECT 214.150 64.845 214.380 65.160 ;
        RECT 214.150 64.660 215.265 64.845 ;
        RECT 214.200 64.625 215.265 64.660 ;
        RECT 214.205 63.540 214.540 64.625 ;
        RECT 215.045 64.510 215.265 64.625 ;
        RECT 216.080 64.510 216.310 64.670 ;
        RECT 215.045 64.290 216.310 64.510 ;
        RECT 216.080 63.670 216.310 64.290 ;
        RECT 213.640 60.240 214.640 63.540 ;
      LAYER via ;
        RECT 213.895 60.465 214.475 61.045 ;
      LAYER met2 ;
        RECT 213.640 0.000 214.640 61.650 ;
        RECT 213.640 -3.280 213.920 0.000 ;
    END
  END dout
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER li1 ;
        RECT 210.985 110.720 211.315 111.210 ;
        RECT 207.150 110.030 207.480 110.520 ;
        RECT 214.830 103.340 216.990 103.690 ;
        RECT 206.680 99.360 206.850 99.860 ;
        RECT 207.650 99.360 207.820 99.860 ;
        RECT 210.750 98.240 210.920 98.740 ;
        RECT 211.810 98.240 211.980 98.740 ;
        RECT 204.020 91.580 204.480 91.750 ;
      LAYER mcon ;
        RECT 211.065 110.880 211.235 111.050 ;
        RECT 207.230 110.190 207.400 110.360 ;
        RECT 214.925 103.430 215.095 103.600 ;
        RECT 215.285 103.430 215.455 103.600 ;
        RECT 215.645 103.430 215.815 103.600 ;
        RECT 216.005 103.430 216.175 103.600 ;
        RECT 216.365 103.430 216.535 103.600 ;
        RECT 216.725 103.430 216.895 103.600 ;
        RECT 206.680 99.525 206.850 99.695 ;
        RECT 207.650 99.525 207.820 99.695 ;
        RECT 210.750 98.405 210.920 98.575 ;
        RECT 211.810 98.405 211.980 98.575 ;
        RECT 204.165 91.580 204.335 91.750 ;
      LAYER met1 ;
        RECT 218.280 116.060 219.280 117.060 ;
        RECT 213.210 115.665 213.535 115.755 ;
        RECT 218.665 115.665 218.840 116.060 ;
        RECT 213.210 115.490 218.840 115.665 ;
        RECT 213.210 114.650 213.535 115.490 ;
        RECT 210.955 111.075 211.345 111.190 ;
        RECT 213.220 111.075 213.545 111.545 ;
        RECT 209.630 110.840 213.545 111.075 ;
        RECT 207.120 110.390 207.510 110.500 ;
        RECT 209.630 110.390 209.865 110.840 ;
        RECT 210.955 110.740 211.345 110.840 ;
        RECT 213.220 110.440 213.545 110.840 ;
        RECT 207.120 110.155 209.865 110.390 ;
        RECT 207.120 110.050 207.510 110.155 ;
        RECT 213.155 103.625 213.480 104.425 ;
        RECT 214.835 103.640 215.215 103.655 ;
        RECT 216.675 103.640 216.925 103.690 ;
        RECT 214.835 103.625 216.965 103.640 ;
        RECT 213.155 103.435 216.965 103.625 ;
        RECT 213.155 103.320 213.480 103.435 ;
        RECT 214.835 103.390 216.965 103.435 ;
        RECT 214.835 103.385 215.215 103.390 ;
        RECT 206.650 99.690 206.880 99.840 ;
        RECT 207.620 99.690 207.850 99.840 ;
        RECT 206.650 99.515 208.430 99.690 ;
        RECT 206.650 99.380 206.880 99.515 ;
        RECT 207.620 99.380 207.850 99.515 ;
        RECT 208.210 99.410 208.430 99.515 ;
        RECT 208.210 98.545 208.535 99.410 ;
        RECT 210.720 98.545 210.950 98.720 ;
        RECT 211.780 98.545 212.010 98.720 ;
        RECT 213.215 98.545 213.540 99.390 ;
        RECT 208.210 98.370 213.540 98.545 ;
        RECT 208.210 98.305 208.535 98.370 ;
        RECT 210.720 98.260 210.950 98.370 ;
        RECT 211.780 98.260 212.010 98.370 ;
        RECT 213.215 98.285 213.540 98.370 ;
        RECT 208.185 92.685 208.510 93.030 ;
        RECT 204.140 92.485 208.510 92.685 ;
        RECT 204.140 91.780 204.340 92.485 ;
        RECT 208.185 91.925 208.510 92.485 ;
        RECT 204.040 91.550 204.460 91.780 ;
      LAYER via ;
        RECT 218.460 116.285 219.040 116.865 ;
        RECT 213.240 115.395 213.500 115.655 ;
        RECT 213.240 115.075 213.500 115.335 ;
        RECT 213.240 114.755 213.500 115.015 ;
        RECT 213.250 111.185 213.510 111.445 ;
        RECT 213.250 110.865 213.510 111.125 ;
        RECT 213.250 110.545 213.510 110.805 ;
        RECT 213.185 104.065 213.445 104.325 ;
        RECT 213.185 103.745 213.445 104.005 ;
        RECT 213.185 103.425 213.445 103.685 ;
        RECT 208.240 99.050 208.500 99.310 ;
        RECT 208.240 98.730 208.500 98.990 ;
        RECT 213.245 99.030 213.505 99.290 ;
        RECT 208.240 98.410 208.500 98.670 ;
        RECT 213.245 98.710 213.505 98.970 ;
        RECT 213.245 98.390 213.505 98.650 ;
        RECT 208.215 92.670 208.475 92.930 ;
        RECT 208.215 92.350 208.475 92.610 ;
        RECT 208.215 92.030 208.475 92.290 ;
      LAYER met2 ;
        RECT 519.780 135.970 520.420 218.525 ;
        RECT 218.280 134.970 520.420 135.970 ;
        RECT 218.280 116.060 219.280 134.970 ;
        RECT 213.160 114.700 213.585 115.705 ;
        RECT 213.285 111.495 213.460 114.700 ;
        RECT 213.170 110.490 213.595 111.495 ;
        RECT 213.285 104.375 213.460 110.490 ;
        RECT 213.105 103.370 213.530 104.375 ;
        RECT 208.160 98.355 208.585 99.360 ;
        RECT 213.285 99.340 213.460 103.370 ;
        RECT 208.255 92.980 208.430 98.355 ;
        RECT 213.165 98.335 213.590 99.340 ;
        RECT 208.135 91.975 208.560 92.980 ;
    END
  END in
  PIN ena
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER li1 ;
        RECT 205.050 72.760 205.220 73.260 ;
        RECT 206.020 72.760 206.190 73.260 ;
        RECT 207.930 64.570 208.100 64.900 ;
        RECT 209.525 64.570 209.695 64.900 ;
      LAYER mcon ;
        RECT 205.050 72.925 205.220 73.095 ;
        RECT 206.020 72.925 206.190 73.095 ;
        RECT 207.930 64.650 208.100 64.820 ;
        RECT 209.525 64.650 209.695 64.820 ;
      LAYER met1 ;
        RECT 205.020 73.080 205.250 73.240 ;
        RECT 205.990 73.080 206.220 73.240 ;
        RECT 207.800 73.080 208.130 73.130 ;
        RECT 205.020 72.880 208.130 73.080 ;
        RECT 205.020 72.780 205.250 72.880 ;
        RECT 205.990 72.780 206.230 72.880 ;
        RECT 207.800 72.540 208.130 72.880 ;
        RECT 207.900 64.810 208.130 64.880 ;
        RECT 208.710 64.810 209.080 64.860 ;
        RECT 209.495 64.810 209.725 64.880 ;
        RECT 207.880 64.570 209.740 64.810 ;
        RECT 208.710 64.390 209.080 64.570 ;
        RECT 208.390 62.540 209.390 64.390 ;
      LAYER via ;
        RECT 207.835 72.705 208.095 72.965 ;
        RECT 208.765 64.480 209.025 64.740 ;
        RECT 208.620 62.815 209.200 63.395 ;
      LAYER met2 ;
        RECT 207.750 72.590 208.180 73.080 ;
        RECT 207.820 65.750 208.090 72.590 ;
        RECT 207.820 65.480 209.025 65.750 ;
        RECT 208.755 64.810 209.025 65.480 ;
        RECT 208.660 64.410 209.130 64.810 ;
        RECT 208.390 0.000 209.390 63.540 ;
        RECT 208.390 -3.280 208.670 0.000 ;
    END
  END ena
  PIN stdby
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER li1 ;
        RECT 224.270 72.760 224.440 73.260 ;
        RECT 225.240 72.760 225.410 73.260 ;
        RECT 220.765 64.570 220.935 64.900 ;
        RECT 222.360 64.570 222.530 64.900 ;
      LAYER mcon ;
        RECT 224.270 72.925 224.440 73.095 ;
        RECT 225.240 72.925 225.410 73.095 ;
        RECT 220.765 64.650 220.935 64.820 ;
        RECT 222.360 64.650 222.530 64.820 ;
      LAYER met1 ;
        RECT 222.330 73.080 222.660 73.130 ;
        RECT 224.240 73.080 224.470 73.240 ;
        RECT 225.210 73.080 225.440 73.240 ;
        RECT 222.330 72.880 225.440 73.080 ;
        RECT 222.330 72.540 222.660 72.880 ;
        RECT 224.230 72.780 224.470 72.880 ;
        RECT 225.210 72.780 225.440 72.880 ;
        RECT 220.735 64.810 220.965 64.880 ;
        RECT 221.380 64.810 221.750 64.860 ;
        RECT 222.330 64.810 222.560 64.880 ;
        RECT 220.720 64.570 222.580 64.810 ;
        RECT 221.380 64.390 221.750 64.570 ;
        RECT 221.070 62.540 222.070 64.390 ;
      LAYER via ;
        RECT 222.365 72.705 222.625 72.965 ;
        RECT 221.435 64.480 221.695 64.740 ;
        RECT 221.270 62.785 221.850 63.365 ;
      LAYER met2 ;
        RECT 222.280 72.590 222.710 73.080 ;
        RECT 222.370 65.750 222.640 72.590 ;
        RECT 221.435 65.480 222.640 65.750 ;
        RECT 221.435 64.810 221.705 65.480 ;
        RECT 221.330 64.410 221.800 64.810 ;
        RECT 221.070 0.000 222.070 63.540 ;
        RECT 221.075 -3.280 221.355 0.000 ;
    END
  END stdby
  PIN out
    PORT
      LAYER li1 ;
        RECT 203.560 113.405 205.720 113.755 ;
      LAYER mcon ;
        RECT 203.655 113.495 203.825 113.665 ;
        RECT 204.015 113.495 204.185 113.665 ;
        RECT 204.375 113.495 204.545 113.665 ;
        RECT 204.735 113.495 204.905 113.665 ;
        RECT 205.095 113.495 205.265 113.665 ;
        RECT 205.455 113.495 205.625 113.665 ;
      LAYER met1 ;
        RECT 209.590 116.060 210.590 117.060 ;
        RECT 210.000 115.295 210.305 116.060 ;
        RECT 205.360 114.990 210.305 115.295 ;
        RECT 205.360 113.705 205.665 114.990 ;
        RECT 203.590 113.455 205.695 113.705 ;
        RECT 205.360 113.420 205.665 113.455 ;
      LAYER via ;
        RECT 209.815 116.290 210.395 116.870 ;
      LAYER met2 ;
        RECT 74.780 135.970 75.420 218.525 ;
        RECT 74.780 134.970 210.590 135.970 ;
        RECT 209.590 116.060 210.590 134.970 ;
    END
  END out
  PIN vssd1
    ANTENNADIFFAREA 21.305099 ;
    PORT
      LAYER pwell ;
        RECT 201.290 66.790 229.085 67.300 ;
        RECT 201.290 62.930 201.800 66.790 ;
        RECT 204.420 64.510 205.150 65.840 ;
        RECT 206.050 63.730 208.740 65.740 ;
        RECT 213.040 63.970 215.050 66.160 ;
        RECT 221.720 63.730 224.410 65.740 ;
        RECT 225.310 64.510 226.040 65.840 ;
        RECT 228.575 62.930 229.085 66.790 ;
        RECT 201.290 62.420 229.085 62.930 ;
      LAYER li1 ;
        RECT 201.420 66.920 228.955 68.055 ;
        RECT 201.420 65.440 208.610 66.920 ;
        RECT 201.420 64.030 206.370 65.440 ;
        RECT 206.720 64.430 207.760 64.600 ;
        RECT 208.440 64.030 208.610 65.440 ;
        RECT 201.420 63.860 208.610 64.030 ;
        RECT 212.810 66.030 213.380 66.920 ;
        RECT 212.810 65.860 214.920 66.030 ;
        RECT 212.810 64.270 213.340 65.860 ;
        RECT 213.740 64.640 213.910 65.180 ;
        RECT 214.750 64.280 214.920 65.860 ;
        RECT 221.855 65.820 228.955 66.920 ;
        RECT 221.850 65.440 228.955 65.820 ;
        RECT 214.750 64.270 214.930 64.280 ;
        RECT 201.420 63.830 206.370 63.860 ;
        RECT 201.420 62.800 206.150 63.830 ;
        RECT 212.810 62.800 214.930 64.270 ;
        RECT 221.850 64.030 222.020 65.440 ;
        RECT 222.700 64.430 223.740 64.600 ;
        RECT 224.090 64.030 228.955 65.440 ;
        RECT 221.850 63.860 228.955 64.030 ;
        RECT 224.090 63.830 228.955 63.860 ;
        RECT 224.185 62.800 228.955 63.830 ;
        RECT 201.420 62.550 228.955 62.800 ;
      LAYER mcon ;
        RECT 201.655 67.315 228.825 67.845 ;
        RECT 201.930 63.740 202.820 66.430 ;
        RECT 205.360 64.630 205.890 65.160 ;
        RECT 206.975 64.430 207.145 64.600 ;
        RECT 207.335 64.430 207.505 64.600 ;
        RECT 213.050 66.525 213.220 66.695 ;
        RECT 213.050 66.165 213.220 66.335 ;
        RECT 213.050 65.805 213.220 65.975 ;
        RECT 213.050 65.445 213.220 65.615 ;
        RECT 213.050 65.085 213.220 65.255 ;
        RECT 213.740 64.825 213.910 64.995 ;
        RECT 224.570 64.630 225.100 65.160 ;
        RECT 222.955 64.430 223.125 64.600 ;
        RECT 223.315 64.430 223.485 64.600 ;
        RECT 227.495 63.270 228.385 66.320 ;
      LAYER met1 ;
        RECT 201.455 66.635 228.980 68.160 ;
        RECT 201.460 64.420 206.280 66.635 ;
        RECT 212.785 65.160 213.705 66.635 ;
        RECT 212.785 64.660 213.940 65.160 ;
        RECT 201.460 64.410 206.340 64.420 ;
        RECT 206.740 64.410 207.740 64.630 ;
        RECT 212.785 64.575 213.810 64.660 ;
        RECT 212.785 64.565 213.705 64.575 ;
        RECT 222.720 64.410 223.720 64.630 ;
        RECT 224.180 64.420 228.980 66.635 ;
        RECT 224.120 64.410 228.980 64.420 ;
        RECT 201.460 64.180 207.750 64.410 ;
        RECT 222.710 64.180 228.980 64.410 ;
        RECT 201.460 63.520 206.280 64.180 ;
        RECT 185.745 62.540 206.280 63.520 ;
        RECT 224.180 62.550 228.980 64.180 ;
      LAYER via ;
        RECT 187.325 62.565 188.865 63.465 ;
        RECT 192.650 62.550 194.190 63.450 ;
      LAYER met2 ;
        RECT 185.745 62.540 196.140 63.520 ;
      LAYER via2 ;
        RECT 187.345 63.100 187.625 63.380 ;
        RECT 187.745 63.100 188.025 63.380 ;
        RECT 188.145 63.100 188.425 63.380 ;
        RECT 188.545 63.100 188.825 63.380 ;
        RECT 192.670 63.100 192.950 63.380 ;
        RECT 193.070 63.100 193.350 63.380 ;
        RECT 193.470 63.100 193.750 63.380 ;
        RECT 193.870 63.100 194.150 63.380 ;
        RECT 187.345 62.655 187.625 62.935 ;
        RECT 187.745 62.655 188.025 62.935 ;
        RECT 188.145 62.655 188.425 62.935 ;
        RECT 188.545 62.655 188.825 62.935 ;
        RECT 192.670 62.630 192.950 62.910 ;
        RECT 193.070 62.630 193.350 62.910 ;
        RECT 193.470 62.630 193.750 62.910 ;
        RECT 193.870 62.630 194.150 62.910 ;
      LAYER met3 ;
        RECT 186.875 62.530 195.000 63.540 ;
      LAYER via3 ;
        RECT 187.325 63.080 187.645 63.400 ;
        RECT 187.725 63.080 188.045 63.400 ;
        RECT 188.125 63.080 188.445 63.400 ;
        RECT 188.525 63.080 188.845 63.400 ;
        RECT 192.650 63.080 192.970 63.400 ;
        RECT 193.050 63.080 193.370 63.400 ;
        RECT 193.450 63.080 193.770 63.400 ;
        RECT 193.850 63.080 194.170 63.400 ;
        RECT 187.325 62.635 187.645 62.955 ;
        RECT 187.725 62.635 188.045 62.955 ;
        RECT 188.125 62.635 188.445 62.955 ;
        RECT 188.525 62.635 188.845 62.955 ;
        RECT 192.650 62.610 192.970 62.930 ;
        RECT 193.050 62.610 193.370 62.930 ;
        RECT 193.450 62.610 193.770 62.930 ;
        RECT 193.850 62.610 194.170 62.930 ;
      LAYER met4 ;
        RECT 187.275 0.000 188.875 211.800 ;
        RECT 192.605 0.000 194.205 211.800 ;
    END
  END vssd1
  PIN vdda1
    ANTENNADIFFAREA 98.890800 ;
    PORT
      LAYER nwell ;
        RECT 201.000 115.450 229.480 117.060 ;
        RECT 201.000 71.320 202.590 115.450 ;
        RECT 206.400 109.360 208.230 111.190 ;
        RECT 209.670 84.630 213.060 109.270 ;
        RECT 207.430 74.510 223.030 77.590 ;
        RECT 207.440 71.320 223.020 74.510 ;
        RECT 227.870 71.320 229.480 115.450 ;
        RECT 201.000 69.710 229.480 71.320 ;
      LAYER li1 ;
        RECT 201.445 115.895 229.015 116.595 ;
        RECT 201.445 70.345 201.615 115.895 ;
        RECT 214.840 114.190 217.000 114.540 ;
        RECT 206.580 110.840 208.050 111.010 ;
        RECT 206.580 109.710 206.750 110.840 ;
        RECT 207.880 109.710 208.050 110.840 ;
        RECT 206.580 109.540 208.050 109.710 ;
        RECT 209.480 108.710 213.270 109.315 ;
        RECT 209.480 106.750 210.250 108.710 ;
        RECT 211.135 108.040 211.595 108.210 ;
        RECT 212.500 106.750 213.270 108.710 ;
        RECT 209.480 106.580 213.270 106.750 ;
        RECT 209.480 105.800 210.250 106.580 ;
        RECT 212.500 105.800 213.270 106.580 ;
        RECT 209.480 105.630 213.270 105.800 ;
        RECT 209.480 103.670 210.250 105.630 ;
        RECT 211.135 104.960 211.595 105.130 ;
        RECT 212.500 103.670 213.270 105.630 ;
        RECT 209.480 103.500 213.270 103.670 ;
        RECT 209.480 102.720 210.250 103.500 ;
        RECT 212.500 102.720 213.270 103.500 ;
        RECT 209.480 102.550 213.270 102.720 ;
        RECT 209.480 100.590 210.250 102.550 ;
        RECT 211.135 101.880 211.595 102.050 ;
        RECT 212.500 100.590 213.270 102.550 ;
        RECT 209.480 100.420 213.270 100.590 ;
        RECT 209.480 99.640 210.250 100.420 ;
        RECT 212.500 99.640 213.270 100.420 ;
        RECT 209.480 99.470 213.270 99.640 ;
        RECT 209.480 97.510 210.250 99.470 ;
        RECT 212.500 97.510 213.270 99.470 ;
        RECT 209.480 97.340 213.270 97.510 ;
        RECT 209.480 96.560 210.250 97.340 ;
        RECT 212.500 96.560 213.270 97.340 ;
        RECT 209.480 96.390 213.270 96.560 ;
        RECT 209.480 94.430 210.250 96.390 ;
        RECT 211.135 95.720 211.595 95.890 ;
        RECT 212.500 94.430 213.270 96.390 ;
        RECT 209.480 94.260 213.270 94.430 ;
        RECT 209.480 93.480 210.250 94.260 ;
        RECT 212.500 93.480 213.270 94.260 ;
        RECT 209.480 93.310 213.270 93.480 ;
        RECT 209.480 91.350 210.250 93.310 ;
        RECT 211.135 92.640 211.595 92.810 ;
        RECT 212.500 91.350 213.270 93.310 ;
        RECT 209.480 91.180 213.270 91.350 ;
        RECT 209.480 90.400 210.250 91.180 ;
        RECT 212.500 90.400 213.270 91.180 ;
        RECT 209.480 90.230 213.270 90.400 ;
        RECT 209.480 88.270 210.250 90.230 ;
        RECT 212.500 88.270 213.270 90.230 ;
        RECT 209.480 88.100 213.270 88.270 ;
        RECT 209.480 87.320 210.250 88.100 ;
        RECT 212.500 87.320 213.270 88.100 ;
        RECT 209.480 87.150 213.270 87.320 ;
        RECT 209.480 85.190 210.250 87.150 ;
        RECT 212.500 85.190 213.270 87.150 ;
        RECT 209.480 85.040 213.270 85.190 ;
        RECT 209.480 85.020 212.670 85.040 ;
        RECT 209.480 85.010 210.250 85.020 ;
        RECT 224.830 80.180 226.990 80.530 ;
        RECT 207.470 76.990 214.220 77.620 ;
        RECT 207.470 75.070 208.010 76.990 ;
        RECT 210.260 75.070 211.340 76.990 ;
        RECT 212.245 75.570 212.705 75.740 ;
        RECT 213.600 75.070 214.220 76.990 ;
        RECT 207.470 73.980 214.220 75.070 ;
        RECT 207.470 72.020 208.010 73.980 ;
        RECT 210.270 73.950 214.220 73.980 ;
        RECT 210.270 72.020 211.340 73.950 ;
        RECT 212.245 73.280 212.705 73.450 ;
        RECT 207.470 72.010 211.340 72.020 ;
        RECT 213.600 72.010 214.220 73.950 ;
        RECT 207.470 71.380 214.220 72.010 ;
        RECT 216.240 76.990 222.990 77.620 ;
        RECT 216.240 75.070 216.860 76.990 ;
        RECT 217.755 75.570 218.215 75.740 ;
        RECT 219.120 75.070 220.200 76.990 ;
        RECT 222.450 75.070 222.990 76.990 ;
        RECT 216.240 73.980 222.990 75.070 ;
        RECT 216.240 73.950 220.190 73.980 ;
        RECT 216.240 72.010 216.860 73.950 ;
        RECT 217.755 73.280 218.215 73.450 ;
        RECT 219.120 72.020 220.190 73.950 ;
        RECT 222.450 72.020 222.990 73.980 ;
        RECT 219.120 72.010 222.990 72.020 ;
        RECT 216.240 71.380 222.990 72.010 ;
        RECT 228.845 70.345 229.015 115.895 ;
        RECT 201.445 69.185 229.015 70.345 ;
      LAYER mcon ;
        RECT 201.755 116.170 201.925 116.340 ;
        RECT 202.115 116.170 202.285 116.340 ;
        RECT 202.475 116.170 202.645 116.340 ;
        RECT 202.835 116.170 203.005 116.340 ;
        RECT 203.195 116.170 203.365 116.340 ;
        RECT 203.555 116.170 203.725 116.340 ;
        RECT 203.915 116.170 204.085 116.340 ;
        RECT 204.275 116.170 204.445 116.340 ;
        RECT 204.635 116.170 204.805 116.340 ;
        RECT 204.995 116.170 205.165 116.340 ;
        RECT 205.355 116.170 205.525 116.340 ;
        RECT 205.715 116.170 205.885 116.340 ;
        RECT 206.075 116.170 206.245 116.340 ;
        RECT 206.435 116.170 206.605 116.340 ;
        RECT 206.795 116.170 206.965 116.340 ;
        RECT 207.155 116.170 207.325 116.340 ;
        RECT 207.515 116.170 207.685 116.340 ;
        RECT 207.875 116.170 208.045 116.340 ;
        RECT 208.235 116.170 208.405 116.340 ;
        RECT 208.595 116.170 208.765 116.340 ;
        RECT 213.975 116.165 214.145 116.335 ;
        RECT 214.335 116.165 214.505 116.335 ;
        RECT 214.695 116.165 214.865 116.335 ;
        RECT 215.055 116.165 215.225 116.335 ;
        RECT 215.415 116.165 215.585 116.335 ;
        RECT 215.775 116.165 215.945 116.335 ;
        RECT 216.135 116.165 216.305 116.335 ;
        RECT 216.495 116.165 216.665 116.335 ;
        RECT 216.855 116.165 217.025 116.335 ;
        RECT 217.215 116.165 217.385 116.335 ;
        RECT 221.310 116.145 221.480 116.315 ;
        RECT 221.670 116.145 221.840 116.315 ;
        RECT 222.030 116.145 222.200 116.315 ;
        RECT 222.390 116.145 222.560 116.315 ;
        RECT 222.750 116.145 222.920 116.315 ;
        RECT 223.110 116.145 223.280 116.315 ;
        RECT 223.470 116.145 223.640 116.315 ;
        RECT 223.830 116.145 224.000 116.315 ;
        RECT 224.190 116.145 224.360 116.315 ;
        RECT 224.550 116.145 224.720 116.315 ;
        RECT 224.910 116.145 225.080 116.315 ;
        RECT 225.270 116.145 225.440 116.315 ;
        RECT 225.630 116.145 225.800 116.315 ;
        RECT 225.990 116.145 226.160 116.315 ;
        RECT 226.350 116.145 226.520 116.315 ;
        RECT 226.710 116.145 226.880 116.315 ;
        RECT 227.070 116.145 227.240 116.315 ;
        RECT 227.430 116.145 227.600 116.315 ;
        RECT 227.790 116.145 227.960 116.315 ;
        RECT 228.150 116.145 228.320 116.315 ;
        RECT 228.510 116.145 228.680 116.315 ;
        RECT 214.935 114.280 215.105 114.450 ;
        RECT 215.295 114.280 215.465 114.450 ;
        RECT 215.655 114.280 215.825 114.450 ;
        RECT 216.015 114.280 216.185 114.450 ;
        RECT 216.375 114.280 216.545 114.450 ;
        RECT 216.735 114.280 216.905 114.450 ;
        RECT 209.605 108.245 210.135 108.775 ;
        RECT 211.280 108.040 211.450 108.210 ;
        RECT 209.610 105.180 210.140 107.150 ;
        RECT 211.280 104.960 211.450 105.130 ;
        RECT 209.600 99.010 210.130 103.500 ;
        RECT 211.280 101.880 211.450 102.050 ;
        RECT 212.630 99.765 213.160 102.815 ;
        RECT 209.595 95.950 210.125 97.560 ;
        RECT 211.280 95.720 211.450 95.890 ;
        RECT 209.595 92.845 210.125 94.455 ;
        RECT 212.655 93.850 213.185 96.900 ;
        RECT 211.280 92.640 211.450 92.810 ;
        RECT 212.630 89.260 213.160 91.230 ;
        RECT 224.920 80.270 225.090 80.440 ;
        RECT 225.280 80.270 225.450 80.440 ;
        RECT 225.640 80.270 225.810 80.440 ;
        RECT 226.000 80.270 226.170 80.440 ;
        RECT 226.360 80.270 226.530 80.440 ;
        RECT 226.720 80.270 226.890 80.440 ;
        RECT 213.110 77.230 213.280 77.400 ;
        RECT 213.470 77.230 213.640 77.400 ;
        RECT 213.830 77.230 214.000 77.400 ;
        RECT 212.390 75.570 212.560 75.740 ;
        RECT 212.440 74.235 214.050 74.765 ;
        RECT 212.390 73.280 212.560 73.450 ;
        RECT 213.165 71.600 213.335 71.770 ;
        RECT 213.525 71.600 213.695 71.770 ;
        RECT 213.885 71.600 214.055 71.770 ;
        RECT 216.460 77.230 216.630 77.400 ;
        RECT 216.820 77.230 216.990 77.400 ;
        RECT 217.180 77.230 217.350 77.400 ;
        RECT 217.900 75.570 218.070 75.740 ;
        RECT 216.410 74.235 218.020 74.765 ;
        RECT 217.900 73.280 218.070 73.450 ;
        RECT 216.405 71.600 216.575 71.770 ;
        RECT 216.765 71.600 216.935 71.770 ;
        RECT 217.125 71.600 217.295 71.770 ;
        RECT 201.655 69.385 228.825 69.915 ;
      LAYER met1 ;
        RECT 201.545 115.970 208.970 116.530 ;
        RECT 213.770 115.960 217.610 116.515 ;
        RECT 221.225 116.465 228.770 116.485 ;
        RECT 221.165 115.990 228.830 116.465 ;
        RECT 221.225 115.970 228.770 115.990 ;
        RECT 214.840 114.190 217.000 115.170 ;
        RECT 209.500 108.890 210.240 108.910 ;
        RECT 209.440 108.545 210.300 108.890 ;
        RECT 209.440 108.140 211.585 108.545 ;
        RECT 209.440 108.130 210.300 108.140 ;
        RECT 209.500 108.110 210.240 108.130 ;
        RECT 211.155 108.010 211.575 108.140 ;
        RECT 209.470 105.455 210.280 107.330 ;
        RECT 209.470 105.050 211.585 105.455 ;
        RECT 209.470 105.000 210.280 105.050 ;
        RECT 211.155 104.930 211.575 105.050 ;
        RECT 209.465 102.375 210.270 103.600 ;
        RECT 212.565 102.950 214.345 102.970 ;
        RECT 209.465 101.970 211.575 102.375 ;
        RECT 209.465 98.910 210.270 101.970 ;
        RECT 211.155 101.850 211.575 101.970 ;
        RECT 212.540 99.630 214.345 102.950 ;
        RECT 212.565 99.625 214.345 99.630 ;
        RECT 209.465 97.240 210.260 97.700 ;
        RECT 213.775 97.240 214.345 99.625 ;
        RECT 209.465 97.090 214.345 97.240 ;
        RECT 209.465 95.860 214.340 97.090 ;
        RECT 209.465 95.855 211.595 95.860 ;
        RECT 209.465 95.805 210.260 95.855 ;
        RECT 211.155 95.690 211.575 95.855 ;
        RECT 209.465 94.430 210.260 94.595 ;
        RECT 212.565 94.430 214.340 95.860 ;
        RECT 209.465 93.445 214.340 94.430 ;
        RECT 209.465 93.110 214.355 93.445 ;
        RECT 209.465 92.730 211.605 93.110 ;
        RECT 209.465 92.700 210.260 92.730 ;
        RECT 211.155 92.610 211.575 92.730 ;
        RECT 212.830 91.340 214.355 93.110 ;
        RECT 212.520 91.215 214.355 91.340 ;
        RECT 212.520 89.205 214.350 91.215 ;
        RECT 212.525 89.185 213.265 89.205 ;
        RECT 224.830 80.175 226.995 82.220 ;
        RECT 212.850 77.000 217.610 77.630 ;
        RECT 212.265 75.740 212.685 75.770 ;
        RECT 212.260 75.480 212.690 75.740 ;
        RECT 213.595 75.480 216.865 77.000 ;
        RECT 217.775 75.740 218.195 75.770 ;
        RECT 217.770 75.480 218.200 75.740 ;
        RECT 212.260 73.590 218.200 75.480 ;
        RECT 212.260 73.270 212.690 73.590 ;
        RECT 212.265 73.250 212.685 73.270 ;
        RECT 213.595 72.000 216.865 73.590 ;
        RECT 217.770 73.270 218.200 73.590 ;
        RECT 217.775 73.250 218.195 73.270 ;
        RECT 213.000 71.370 217.460 72.000 ;
        RECT 213.000 70.765 216.385 71.370 ;
        RECT 201.420 68.975 229.045 70.765 ;
      LAYER via ;
        RECT 221.345 116.100 221.605 116.360 ;
        RECT 221.665 116.100 221.925 116.360 ;
        RECT 221.985 116.100 222.245 116.360 ;
        RECT 222.305 116.100 222.565 116.360 ;
        RECT 222.625 116.100 222.885 116.360 ;
        RECT 222.945 116.100 223.205 116.360 ;
        RECT 223.265 116.100 223.525 116.360 ;
        RECT 223.585 116.100 223.845 116.360 ;
        RECT 223.905 116.100 224.165 116.360 ;
        RECT 224.225 116.100 224.485 116.360 ;
        RECT 224.545 116.100 224.805 116.360 ;
        RECT 224.865 116.100 225.125 116.360 ;
        RECT 225.185 116.100 225.445 116.360 ;
        RECT 225.505 116.100 225.765 116.360 ;
        RECT 225.825 116.100 226.085 116.360 ;
        RECT 226.145 116.100 226.405 116.360 ;
        RECT 226.465 116.100 226.725 116.360 ;
        RECT 226.785 116.100 227.045 116.360 ;
        RECT 227.105 116.100 227.365 116.360 ;
        RECT 227.425 116.100 227.685 116.360 ;
        RECT 227.745 116.100 228.005 116.360 ;
        RECT 228.065 116.100 228.325 116.360 ;
        RECT 228.385 116.100 228.645 116.360 ;
        RECT 214.995 114.405 216.855 114.985 ;
        RECT 209.580 108.220 210.160 108.800 ;
        RECT 209.585 105.075 210.165 107.255 ;
        RECT 209.575 99.045 210.155 103.465 ;
        RECT 209.570 95.985 210.150 97.525 ;
        RECT 209.570 92.880 210.150 94.420 ;
        RECT 213.025 93.285 214.245 97.065 ;
        RECT 213.065 89.455 214.285 91.955 ;
        RECT 224.975 81.380 226.835 81.960 ;
        RECT 224.255 69.095 228.995 70.635 ;
      LAYER met2 ;
        RECT 221.135 115.350 229.275 117.060 ;
        RECT 214.670 114.080 229.275 115.350 ;
        RECT 209.005 92.565 210.860 109.545 ;
        RECT 221.135 97.230 229.275 114.080 ;
        RECT 212.920 93.090 229.275 97.230 ;
        RECT 219.265 93.080 229.275 93.090 ;
        RECT 221.135 92.260 229.275 93.080 ;
        RECT 219.265 92.250 229.275 92.260 ;
        RECT 212.950 89.195 229.275 92.250 ;
        RECT 221.135 83.655 229.275 89.195 ;
        RECT 224.085 79.715 229.275 83.655 ;
        RECT 224.085 68.985 229.285 79.715 ;
      LAYER via2 ;
        RECT 222.435 116.620 222.715 116.900 ;
        RECT 222.835 116.620 223.115 116.900 ;
        RECT 223.235 116.620 223.515 116.900 ;
        RECT 223.635 116.620 223.915 116.900 ;
        RECT 226.580 116.620 226.860 116.900 ;
        RECT 226.980 116.620 227.260 116.900 ;
        RECT 227.380 116.620 227.660 116.900 ;
        RECT 227.780 116.620 228.060 116.900 ;
      LAYER met3 ;
        RECT 221.135 116.435 229.275 117.060 ;
      LAYER via3 ;
        RECT 222.415 116.600 222.735 116.920 ;
        RECT 222.815 116.600 223.135 116.920 ;
        RECT 223.215 116.600 223.535 116.920 ;
        RECT 223.615 116.600 223.935 116.920 ;
        RECT 226.560 116.600 226.880 116.920 ;
        RECT 226.960 116.600 227.280 116.920 ;
        RECT 227.360 116.600 227.680 116.920 ;
        RECT 227.760 116.600 228.080 116.920 ;
      LAYER met4 ;
        RECT 222.405 0.000 224.005 211.800 ;
        RECT 226.550 0.000 228.150 211.800 ;
    END
  END vdda1
  PIN vccd1
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER nwell ;
        RECT 208.830 63.680 211.670 65.790 ;
        RECT 215.360 62.930 217.470 65.770 ;
        RECT 218.790 63.680 221.630 65.790 ;
      LAYER li1 ;
        RECT 211.135 89.560 211.595 89.730 ;
        RECT 209.010 65.440 211.850 65.830 ;
        RECT 209.010 64.030 209.180 65.440 ;
        RECT 211.320 65.100 211.850 65.440 ;
        RECT 215.535 65.410 217.630 66.085 ;
        RECT 209.910 64.430 210.950 64.600 ;
        RECT 211.320 64.310 212.310 65.100 ;
        RECT 211.320 64.030 211.850 64.310 ;
        RECT 209.010 63.860 211.850 64.030 ;
        RECT 211.340 63.840 211.850 63.860 ;
        RECT 215.540 63.280 215.710 65.410 ;
        RECT 216.550 63.650 216.720 64.690 ;
        RECT 217.120 63.280 217.630 65.410 ;
        RECT 218.610 65.440 221.450 65.830 ;
        RECT 218.610 65.100 219.140 65.440 ;
        RECT 218.150 64.310 219.140 65.100 ;
        RECT 219.510 64.430 220.550 64.600 ;
        RECT 218.610 64.030 219.140 64.310 ;
        RECT 221.280 64.030 221.450 65.440 ;
        RECT 218.610 63.860 221.450 64.030 ;
        RECT 218.610 63.840 219.120 63.860 ;
        RECT 215.540 63.110 217.630 63.280 ;
      LAYER mcon ;
        RECT 211.280 89.560 211.450 89.730 ;
        RECT 210.165 64.430 210.335 64.600 ;
        RECT 210.525 64.430 210.695 64.600 ;
        RECT 211.640 64.460 212.170 64.990 ;
        RECT 216.550 64.265 216.720 64.435 ;
        RECT 216.550 63.905 216.720 64.075 ;
        RECT 217.310 64.270 217.480 64.440 ;
        RECT 218.290 64.460 218.820 64.990 ;
        RECT 219.765 64.430 219.935 64.600 ;
        RECT 220.125 64.430 220.295 64.600 ;
        RECT 217.310 63.910 217.480 64.080 ;
      LAYER met1 ;
        RECT 211.140 89.485 211.605 90.795 ;
        RECT 211.315 65.780 212.305 65.785 ;
        RECT 209.930 64.460 210.930 64.630 ;
        RECT 211.310 64.460 212.310 65.780 ;
        RECT 209.930 64.230 212.310 64.460 ;
        RECT 211.310 63.390 212.310 64.230 ;
        RECT 216.520 64.665 216.750 64.670 ;
        RECT 218.150 64.665 219.150 65.800 ;
        RECT 216.520 64.460 219.150 64.665 ;
        RECT 219.530 64.460 220.530 64.630 ;
        RECT 216.520 64.230 220.530 64.460 ;
        RECT 216.520 63.670 219.150 64.230 ;
        RECT 216.670 63.650 219.150 63.670 ;
        RECT 211.315 63.375 212.305 63.390 ;
        RECT 218.150 62.430 219.150 63.650 ;
      LAYER via ;
        RECT 211.240 90.330 211.500 90.590 ;
        RECT 211.240 90.010 211.500 90.270 ;
        RECT 211.240 89.690 211.500 89.950 ;
        RECT 211.515 63.485 212.095 65.665 ;
        RECT 218.205 63.505 219.105 65.685 ;
      LAYER met2 ;
        RECT 208.890 89.515 211.655 90.745 ;
        RECT 208.890 85.410 209.705 89.515 ;
        RECT 208.890 84.430 212.930 85.410 ;
        RECT 212.155 65.785 212.930 84.430 ;
        RECT 211.315 64.920 212.930 65.785 ;
        RECT 218.150 64.920 219.150 65.800 ;
        RECT 211.315 63.380 219.150 64.920 ;
        RECT 211.315 63.375 212.305 63.380 ;
        RECT 215.290 62.430 219.150 63.380 ;
      LAYER via2 ;
        RECT 216.700 62.990 216.980 63.270 ;
        RECT 217.100 62.990 217.380 63.270 ;
        RECT 217.500 62.990 217.780 63.270 ;
        RECT 217.900 62.990 218.180 63.270 ;
        RECT 216.700 62.545 216.980 62.825 ;
        RECT 217.100 62.545 217.380 62.825 ;
        RECT 217.500 62.545 217.780 62.825 ;
        RECT 217.900 62.545 218.180 62.825 ;
      LAYER met3 ;
        RECT 216.230 62.420 219.150 63.430 ;
      LAYER via3 ;
        RECT 216.680 62.970 217.000 63.290 ;
        RECT 217.080 62.970 217.400 63.290 ;
        RECT 217.480 62.970 217.800 63.290 ;
        RECT 217.880 62.970 218.200 63.290 ;
        RECT 216.680 62.525 217.000 62.845 ;
        RECT 217.080 62.525 217.400 62.845 ;
        RECT 217.480 62.525 217.800 62.845 ;
        RECT 217.880 62.525 218.200 62.845 ;
      LAYER met4 ;
        RECT 216.610 0.000 218.210 211.800 ;
    END
  END vccd1
  PIN vssa1
    ANTENNADIFFAREA 81.684601 ;
    PORT
      LAYER pwell ;
        RECT 214.060 114.890 227.780 115.320 ;
        RECT 202.780 114.105 213.500 114.535 ;
        RECT 202.780 113.055 203.210 114.105 ;
        RECT 213.070 113.055 213.500 114.105 ;
        RECT 202.780 112.625 213.500 113.055 ;
        RECT 205.760 111.400 208.870 111.830 ;
        RECT 205.760 109.150 206.190 111.400 ;
        RECT 208.440 109.150 208.870 111.400 ;
        RECT 210.285 110.100 212.015 111.830 ;
        RECT 205.760 108.720 208.870 109.150 ;
        RECT 202.800 103.830 205.700 106.510 ;
        RECT 205.800 103.830 208.700 106.510 ;
        RECT 214.060 106.370 214.490 114.890 ;
        RECT 227.350 106.370 227.780 114.890 ;
        RECT 214.060 105.940 227.780 106.370 ;
        RECT 214.050 104.040 227.770 104.470 ;
        RECT 202.800 101.050 205.700 103.730 ;
        RECT 205.800 101.050 208.700 103.730 ;
        RECT 202.800 98.270 205.700 100.950 ;
        RECT 205.800 98.270 208.700 100.950 ;
        RECT 202.800 95.490 205.700 98.170 ;
        RECT 202.800 92.710 205.700 95.390 ;
        RECT 205.800 92.710 208.700 95.390 ;
        RECT 202.800 89.930 205.700 92.610 ;
        RECT 205.800 89.930 208.700 92.610 ;
        RECT 202.800 87.150 205.700 89.830 ;
        RECT 205.800 87.150 208.700 89.830 ;
        RECT 202.765 83.895 213.485 84.325 ;
        RECT 202.765 82.015 203.195 83.895 ;
        RECT 213.055 82.015 213.485 83.895 ;
        RECT 214.050 83.070 214.480 104.040 ;
        RECT 227.340 83.070 227.770 104.040 ;
        RECT 214.050 82.640 227.770 83.070 ;
        RECT 202.765 81.585 213.485 82.015 ;
        RECT 212.050 80.880 227.770 81.310 ;
        RECT 212.050 79.830 212.480 80.880 ;
        RECT 227.340 79.830 227.770 80.880 ;
        RECT 212.050 79.400 227.770 79.830 ;
        RECT 204.180 74.700 207.080 77.380 ;
        RECT 223.380 74.700 226.280 77.380 ;
        RECT 204.170 71.670 207.070 74.350 ;
        RECT 223.390 71.670 226.290 74.350 ;
      LAYER li1 ;
        RECT 213.285 115.190 214.340 115.200 ;
        RECT 227.460 115.190 228.200 115.210 ;
        RECT 213.285 115.020 228.200 115.190 ;
        RECT 213.285 114.405 214.360 115.020 ;
        RECT 202.910 114.235 214.360 114.405 ;
        RECT 202.910 112.925 203.080 114.235 ;
        RECT 213.200 112.925 214.360 114.235 ;
        RECT 202.910 112.860 214.360 112.925 ;
        RECT 202.900 111.615 214.360 112.860 ;
        RECT 205.890 111.530 212.345 111.615 ;
        RECT 205.890 109.020 206.060 111.530 ;
        RECT 208.570 110.400 210.585 111.530 ;
        RECT 211.715 110.400 212.345 111.530 ;
        RECT 208.570 109.865 212.345 110.400 ;
        RECT 208.570 109.020 208.740 109.865 ;
        RECT 205.890 108.850 208.740 109.020 ;
        RECT 202.380 106.145 209.120 106.635 ;
        RECT 202.380 104.190 203.180 106.145 ;
        RECT 204.020 105.480 204.480 105.650 ;
        RECT 205.340 104.190 206.170 106.145 ;
        RECT 208.320 104.190 209.120 106.145 ;
        RECT 202.380 104.020 209.120 104.190 ;
        RECT 202.380 103.540 203.180 104.020 ;
        RECT 205.370 103.540 206.170 104.020 ;
        RECT 208.320 103.540 209.120 104.020 ;
        RECT 202.380 103.370 209.120 103.540 ;
        RECT 202.380 101.410 203.180 103.370 ;
        RECT 204.020 102.700 204.480 102.870 ;
        RECT 205.340 101.410 206.170 103.370 ;
        RECT 208.320 101.410 209.120 103.370 ;
        RECT 202.380 101.240 209.120 101.410 ;
        RECT 202.380 100.760 203.180 101.240 ;
        RECT 205.370 100.760 206.170 101.240 ;
        RECT 208.320 100.760 209.120 101.240 ;
        RECT 202.380 100.590 209.120 100.760 ;
        RECT 202.380 98.630 203.180 100.590 ;
        RECT 204.020 99.920 204.480 100.090 ;
        RECT 205.340 98.630 206.170 100.590 ;
        RECT 208.320 98.630 209.120 100.590 ;
        RECT 202.380 98.460 209.120 98.630 ;
        RECT 202.380 97.980 203.180 98.460 ;
        RECT 205.370 97.980 206.170 98.460 ;
        RECT 202.380 97.810 206.170 97.980 ;
        RECT 202.380 95.850 203.180 97.810 ;
        RECT 204.020 96.350 204.480 96.520 ;
        RECT 205.340 95.850 206.170 97.810 ;
        RECT 202.380 95.680 206.170 95.850 ;
        RECT 202.380 95.200 203.180 95.680 ;
        RECT 205.370 95.200 206.170 95.680 ;
        RECT 208.320 95.200 209.120 98.460 ;
        RECT 202.380 95.030 209.120 95.200 ;
        RECT 202.380 93.070 203.180 95.030 ;
        RECT 204.020 94.360 204.480 94.530 ;
        RECT 205.340 93.070 206.170 95.030 ;
        RECT 207.020 94.360 207.480 94.530 ;
        RECT 208.320 93.070 209.120 95.030 ;
        RECT 202.380 92.900 209.120 93.070 ;
        RECT 202.380 92.420 203.180 92.900 ;
        RECT 205.370 92.420 206.170 92.900 ;
        RECT 208.320 92.420 209.120 92.900 ;
        RECT 202.380 92.250 209.120 92.420 ;
        RECT 202.380 90.290 203.180 92.250 ;
        RECT 205.340 90.290 206.170 92.250 ;
        RECT 207.020 91.580 207.480 91.750 ;
        RECT 208.320 90.290 209.120 92.250 ;
        RECT 202.380 90.120 209.120 90.290 ;
        RECT 202.380 89.640 203.180 90.120 ;
        RECT 205.370 89.640 206.170 90.120 ;
        RECT 208.320 89.640 209.120 90.120 ;
        RECT 202.380 89.470 209.120 89.640 ;
        RECT 202.380 87.510 203.180 89.470 ;
        RECT 205.340 87.510 206.170 89.470 ;
        RECT 207.020 88.800 207.480 88.970 ;
        RECT 208.320 87.510 209.120 89.470 ;
        RECT 202.380 87.360 209.120 87.510 ;
        RECT 202.990 87.340 209.120 87.360 ;
        RECT 205.370 87.320 206.170 87.340 ;
        RECT 208.320 87.330 209.120 87.340 ;
        RECT 213.630 106.240 214.360 111.615 ;
        RECT 227.460 106.240 228.200 115.020 ;
        RECT 213.630 104.170 228.200 106.240 ;
        RECT 213.630 104.075 214.360 104.170 ;
        RECT 213.630 84.570 214.350 104.075 ;
        RECT 227.460 93.860 228.200 104.170 ;
        RECT 227.470 91.635 228.200 93.860 ;
        RECT 202.260 84.025 214.350 84.570 ;
        RECT 202.260 81.885 203.065 84.025 ;
        RECT 213.185 82.940 214.350 84.025 ;
        RECT 227.460 82.940 228.200 91.635 ;
        RECT 210.545 82.365 212.705 82.715 ;
        RECT 213.185 82.170 228.200 82.940 ;
        RECT 213.185 81.885 214.340 82.170 ;
        RECT 202.260 81.880 214.340 81.885 ;
        RECT 202.020 81.740 214.340 81.880 ;
        RECT 227.460 81.740 228.200 82.170 ;
        RECT 202.020 81.015 228.200 81.740 ;
        RECT 202.020 79.485 203.830 81.015 ;
        RECT 205.315 80.520 207.305 81.015 ;
        RECT 211.585 81.010 228.200 81.015 ;
        RECT 211.585 79.700 212.350 81.010 ;
        RECT 227.460 79.700 228.200 81.010 ;
        RECT 211.585 79.130 228.200 79.700 ;
        RECT 227.460 79.110 228.200 79.130 ;
        RECT 203.730 77.000 207.220 77.630 ;
        RECT 203.730 75.070 204.560 77.000 ;
        RECT 205.400 76.350 205.860 76.520 ;
        RECT 206.690 75.070 207.220 77.000 ;
        RECT 203.730 73.990 207.220 75.070 ;
        RECT 203.730 72.050 204.560 73.990 ;
        RECT 205.390 72.530 205.850 72.700 ;
        RECT 206.690 72.050 207.220 73.990 ;
        RECT 203.730 71.420 207.220 72.050 ;
        RECT 223.240 77.000 226.730 77.630 ;
        RECT 223.240 75.070 223.770 77.000 ;
        RECT 224.600 76.350 225.060 76.520 ;
        RECT 225.900 75.070 226.730 77.000 ;
        RECT 223.240 73.990 226.730 75.070 ;
        RECT 223.240 72.050 223.770 73.990 ;
        RECT 224.610 72.530 225.070 72.700 ;
        RECT 225.900 72.050 226.730 73.990 ;
        RECT 223.240 71.420 226.730 72.050 ;
      LAYER mcon ;
        RECT 203.260 111.955 212.790 112.485 ;
        RECT 202.515 87.610 203.045 106.140 ;
        RECT 204.165 105.480 204.335 105.650 ;
        RECT 205.480 105.625 206.010 106.155 ;
        RECT 204.165 102.700 204.335 102.870 ;
        RECT 205.480 102.735 206.010 103.265 ;
        RECT 204.165 99.920 204.335 100.090 ;
        RECT 205.470 99.930 206.000 100.460 ;
        RECT 204.165 96.350 204.335 96.520 ;
        RECT 205.480 94.555 206.010 95.085 ;
        RECT 204.165 94.360 204.335 94.530 ;
        RECT 207.165 94.360 207.335 94.530 ;
        RECT 205.485 88.090 206.015 91.860 ;
        RECT 207.165 91.580 207.335 91.750 ;
        RECT 207.165 88.800 207.335 88.970 ;
        RECT 227.885 114.675 228.055 114.845 ;
        RECT 227.885 114.315 228.055 114.485 ;
        RECT 227.885 113.955 228.055 114.125 ;
        RECT 227.885 113.595 228.055 113.765 ;
        RECT 227.885 113.235 228.055 113.405 ;
        RECT 227.885 112.875 228.055 113.045 ;
        RECT 227.885 112.515 228.055 112.685 ;
        RECT 227.885 112.155 228.055 112.325 ;
        RECT 227.885 111.795 228.055 111.965 ;
        RECT 227.885 111.435 228.055 111.605 ;
        RECT 227.885 111.075 228.055 111.245 ;
        RECT 227.885 110.715 228.055 110.885 ;
        RECT 227.885 110.355 228.055 110.525 ;
        RECT 227.885 109.995 228.055 110.165 ;
        RECT 227.885 109.635 228.055 109.805 ;
        RECT 227.885 109.275 228.055 109.445 ;
        RECT 227.885 108.915 228.055 109.085 ;
        RECT 227.885 108.555 228.055 108.725 ;
        RECT 227.885 108.195 228.055 108.365 ;
        RECT 227.885 107.835 228.055 108.005 ;
        RECT 227.885 107.475 228.055 107.645 ;
        RECT 227.885 107.115 228.055 107.285 ;
        RECT 227.885 106.755 228.055 106.925 ;
        RECT 227.885 106.395 228.055 106.565 ;
        RECT 227.885 106.035 228.055 106.205 ;
        RECT 213.905 104.740 227.395 105.630 ;
        RECT 227.870 103.855 228.040 104.025 ;
        RECT 227.870 103.495 228.040 103.665 ;
        RECT 227.870 103.135 228.040 103.305 ;
        RECT 227.870 102.775 228.040 102.945 ;
        RECT 227.870 102.415 228.040 102.585 ;
        RECT 227.870 102.055 228.040 102.225 ;
        RECT 227.870 101.695 228.040 101.865 ;
        RECT 227.870 101.335 228.040 101.505 ;
        RECT 227.870 100.975 228.040 101.145 ;
        RECT 227.870 100.615 228.040 100.785 ;
        RECT 227.870 100.255 228.040 100.425 ;
        RECT 227.870 99.895 228.040 100.065 ;
        RECT 227.870 99.535 228.040 99.705 ;
        RECT 227.870 99.175 228.040 99.345 ;
        RECT 227.870 98.815 228.040 98.985 ;
        RECT 227.870 98.455 228.040 98.625 ;
        RECT 227.870 98.095 228.040 98.265 ;
        RECT 227.870 97.735 228.040 97.905 ;
        RECT 227.870 97.375 228.040 97.545 ;
        RECT 227.870 97.015 228.040 97.185 ;
        RECT 227.870 96.655 228.040 96.825 ;
        RECT 227.870 96.295 228.040 96.465 ;
        RECT 227.870 95.935 228.040 96.105 ;
        RECT 227.870 95.575 228.040 95.745 ;
        RECT 227.870 95.215 228.040 95.385 ;
        RECT 227.870 94.855 228.040 95.025 ;
        RECT 227.870 94.495 228.040 94.665 ;
        RECT 227.870 94.135 228.040 94.305 ;
        RECT 227.870 93.775 228.040 93.945 ;
        RECT 227.870 93.415 228.040 93.585 ;
        RECT 227.870 93.055 228.040 93.225 ;
        RECT 227.870 92.695 228.040 92.865 ;
        RECT 227.870 92.335 228.040 92.505 ;
        RECT 227.870 91.975 228.040 92.145 ;
        RECT 227.870 91.615 228.040 91.785 ;
        RECT 227.870 91.255 228.040 91.425 ;
        RECT 227.870 90.895 228.040 91.065 ;
        RECT 227.870 90.535 228.040 90.705 ;
        RECT 227.870 90.175 228.040 90.345 ;
        RECT 227.870 89.815 228.040 89.985 ;
        RECT 227.870 89.455 228.040 89.625 ;
        RECT 227.870 89.095 228.040 89.265 ;
        RECT 227.870 88.735 228.040 88.905 ;
        RECT 227.870 88.375 228.040 88.545 ;
        RECT 227.870 88.015 228.040 88.185 ;
        RECT 227.870 87.655 228.040 87.825 ;
        RECT 227.870 87.295 228.040 87.465 ;
        RECT 227.870 86.935 228.040 87.105 ;
        RECT 227.870 86.575 228.040 86.745 ;
        RECT 227.870 86.215 228.040 86.385 ;
        RECT 227.870 85.855 228.040 86.025 ;
        RECT 227.870 85.495 228.040 85.665 ;
        RECT 227.870 85.135 228.040 85.305 ;
        RECT 227.870 84.775 228.040 84.945 ;
        RECT 227.870 84.415 228.040 84.585 ;
        RECT 227.870 84.055 228.040 84.225 ;
        RECT 227.870 83.695 228.040 83.865 ;
        RECT 227.870 83.335 228.040 83.505 ;
        RECT 227.870 82.975 228.040 83.145 ;
        RECT 210.635 82.455 210.805 82.625 ;
        RECT 210.995 82.455 211.165 82.625 ;
        RECT 211.355 82.455 211.525 82.625 ;
        RECT 211.715 82.455 211.885 82.625 ;
        RECT 212.075 82.455 212.245 82.625 ;
        RECT 212.435 82.455 212.605 82.625 ;
        RECT 227.870 82.615 228.040 82.785 ;
        RECT 214.475 82.440 214.645 82.610 ;
        RECT 214.835 82.440 215.005 82.610 ;
        RECT 215.195 82.440 215.365 82.610 ;
        RECT 215.555 82.440 215.725 82.610 ;
        RECT 215.915 82.440 216.085 82.610 ;
        RECT 216.275 82.440 216.445 82.610 ;
        RECT 216.635 82.440 216.805 82.610 ;
        RECT 216.995 82.440 217.165 82.610 ;
        RECT 217.355 82.440 217.525 82.610 ;
        RECT 217.715 82.440 217.885 82.610 ;
        RECT 218.075 82.440 218.245 82.610 ;
        RECT 218.435 82.440 218.605 82.610 ;
        RECT 218.795 82.440 218.965 82.610 ;
        RECT 219.155 82.440 219.325 82.610 ;
        RECT 219.515 82.440 219.685 82.610 ;
        RECT 219.875 82.440 220.045 82.610 ;
        RECT 220.235 82.440 220.405 82.610 ;
        RECT 220.595 82.440 220.765 82.610 ;
        RECT 220.955 82.440 221.125 82.610 ;
        RECT 221.315 82.440 221.485 82.610 ;
        RECT 221.675 82.440 221.845 82.610 ;
        RECT 222.035 82.440 222.205 82.610 ;
        RECT 227.870 82.255 228.040 82.425 ;
        RECT 202.120 79.695 203.730 81.665 ;
        RECT 205.500 80.585 207.110 81.835 ;
        RECT 227.870 81.895 228.040 82.065 ;
        RECT 210.650 81.515 210.820 81.685 ;
        RECT 211.010 81.515 211.180 81.685 ;
        RECT 211.370 81.515 211.540 81.685 ;
        RECT 211.730 81.515 211.900 81.685 ;
        RECT 212.090 81.515 212.260 81.685 ;
        RECT 212.450 81.515 212.620 81.685 ;
        RECT 227.870 81.535 228.040 81.705 ;
        RECT 214.480 81.325 214.650 81.495 ;
        RECT 214.840 81.325 215.010 81.495 ;
        RECT 215.200 81.325 215.370 81.495 ;
        RECT 215.560 81.325 215.730 81.495 ;
        RECT 215.920 81.325 216.090 81.495 ;
        RECT 216.280 81.325 216.450 81.495 ;
        RECT 216.640 81.325 216.810 81.495 ;
        RECT 217.000 81.325 217.170 81.495 ;
        RECT 217.360 81.325 217.530 81.495 ;
        RECT 217.720 81.325 217.890 81.495 ;
        RECT 218.080 81.325 218.250 81.495 ;
        RECT 218.440 81.325 218.610 81.495 ;
        RECT 218.800 81.325 218.970 81.495 ;
        RECT 219.160 81.325 219.330 81.495 ;
        RECT 219.520 81.325 219.690 81.495 ;
        RECT 219.880 81.325 220.050 81.495 ;
        RECT 220.240 81.325 220.410 81.495 ;
        RECT 220.600 81.325 220.770 81.495 ;
        RECT 220.960 81.325 221.130 81.495 ;
        RECT 221.320 81.325 221.490 81.495 ;
        RECT 221.680 81.325 221.850 81.495 ;
        RECT 222.040 81.325 222.210 81.495 ;
        RECT 222.400 81.325 222.570 81.495 ;
        RECT 222.760 81.325 222.930 81.495 ;
        RECT 223.120 81.325 223.290 81.495 ;
        RECT 223.480 81.325 223.650 81.495 ;
        RECT 223.840 81.325 224.010 81.495 ;
        RECT 224.200 81.325 224.370 81.495 ;
        RECT 227.870 81.175 228.040 81.345 ;
        RECT 227.870 80.815 228.040 80.985 ;
        RECT 227.870 80.455 228.040 80.625 ;
        RECT 227.870 80.095 228.040 80.265 ;
        RECT 227.870 79.735 228.040 79.905 ;
        RECT 203.935 76.555 204.105 76.725 ;
        RECT 203.935 76.195 204.105 76.365 ;
        RECT 205.545 76.350 205.715 76.520 ;
        RECT 203.935 75.835 204.105 76.005 ;
        RECT 203.935 75.475 204.105 75.645 ;
        RECT 204.020 74.085 204.910 74.975 ;
        RECT 203.925 73.375 204.095 73.545 ;
        RECT 203.925 73.015 204.095 73.185 ;
        RECT 203.925 72.655 204.095 72.825 ;
        RECT 205.535 72.530 205.705 72.700 ;
        RECT 203.925 72.295 204.095 72.465 ;
        RECT 226.355 76.555 226.525 76.725 ;
        RECT 224.745 76.350 224.915 76.520 ;
        RECT 226.355 76.195 226.525 76.365 ;
        RECT 226.355 75.835 226.525 76.005 ;
        RECT 226.355 75.475 226.525 75.645 ;
        RECT 225.550 74.085 226.440 74.975 ;
        RECT 226.365 73.375 226.535 73.545 ;
        RECT 226.365 73.015 226.535 73.185 ;
        RECT 224.755 72.530 224.925 72.700 ;
        RECT 226.365 72.655 226.535 72.825 ;
        RECT 226.365 72.295 226.535 72.465 ;
      LAYER met1 ;
        RECT 203.040 111.895 213.010 112.570 ;
        RECT 202.380 96.395 203.175 106.370 ;
        RECT 205.370 105.880 206.120 106.315 ;
        RECT 227.470 105.890 228.195 115.355 ;
        RECT 204.040 105.580 206.120 105.880 ;
        RECT 204.040 105.450 204.460 105.580 ;
        RECT 205.370 105.460 206.120 105.580 ;
        RECT 213.725 104.445 228.195 105.890 ;
        RECT 205.370 103.140 206.120 103.425 ;
        RECT 204.050 102.900 206.120 103.140 ;
        RECT 204.040 102.840 206.120 102.900 ;
        RECT 204.040 102.670 204.460 102.840 ;
        RECT 205.370 102.570 206.120 102.840 ;
        RECT 205.360 100.320 206.110 100.620 ;
        RECT 204.040 100.020 206.110 100.320 ;
        RECT 204.040 99.890 204.460 100.020 ;
        RECT 205.360 99.765 206.110 100.020 ;
        RECT 204.040 96.395 204.460 96.550 ;
        RECT 202.380 96.035 204.490 96.395 ;
        RECT 202.380 94.860 203.175 96.035 ;
        RECT 202.380 94.560 204.450 94.860 ;
        RECT 205.370 94.825 206.120 95.245 ;
        RECT 202.380 94.445 204.460 94.560 ;
        RECT 202.380 90.825 203.175 94.445 ;
        RECT 204.040 94.330 204.460 94.445 ;
        RECT 205.350 94.440 207.470 94.825 ;
        RECT 205.370 94.390 206.120 94.440 ;
        RECT 207.040 94.330 207.460 94.440 ;
        RECT 205.375 92.030 206.125 92.090 ;
        RECT 205.370 91.645 207.490 92.030 ;
        RECT 202.380 90.410 203.180 90.825 ;
        RECT 202.380 89.300 203.175 90.410 ;
        RECT 205.375 89.310 206.125 91.645 ;
        RECT 207.040 91.550 207.460 91.645 ;
        RECT 202.380 88.885 203.180 89.300 ;
        RECT 205.375 88.925 207.495 89.310 ;
        RECT 202.380 87.355 203.175 88.885 ;
        RECT 205.375 87.855 206.125 88.925 ;
        RECT 207.040 88.770 207.460 88.925 ;
        RECT 210.545 81.885 212.710 82.715 ;
        RECT 214.320 82.280 222.360 82.760 ;
        RECT 202.020 76.840 203.830 81.880 ;
        RECT 205.315 80.520 207.305 81.885 ;
        RECT 210.535 81.315 212.735 81.885 ;
        RECT 214.335 81.605 224.475 81.650 ;
        RECT 210.545 81.310 212.710 81.315 ;
        RECT 214.335 81.210 224.480 81.605 ;
        RECT 214.335 81.170 224.475 81.210 ;
        RECT 227.470 78.765 228.195 104.445 ;
        RECT 226.870 76.840 228.195 78.765 ;
        RECT 202.020 76.420 205.850 76.840 ;
        RECT 224.610 76.420 228.195 76.840 ;
        RECT 202.020 75.310 204.680 76.420 ;
        RECT 205.420 76.320 205.840 76.420 ;
        RECT 224.620 76.320 225.040 76.420 ;
        RECT 225.780 75.310 228.195 76.420 ;
        RECT 202.020 73.760 205.050 75.310 ;
        RECT 225.410 73.760 228.195 75.310 ;
        RECT 202.020 72.600 204.680 73.760 ;
        RECT 205.410 72.600 205.830 72.730 ;
        RECT 224.630 72.600 225.050 72.730 ;
        RECT 225.780 72.600 228.195 73.760 ;
        RECT 202.020 72.180 205.840 72.600 ;
        RECT 224.620 72.180 228.195 72.600 ;
        RECT 202.020 70.940 203.830 72.180 ;
        RECT 226.870 71.325 228.195 72.180 ;
        RECT 227.470 71.320 228.195 71.325 ;
      LAYER via ;
        RECT 203.130 112.095 203.390 112.355 ;
        RECT 203.450 112.095 203.710 112.355 ;
        RECT 203.770 112.095 204.030 112.355 ;
        RECT 204.090 112.095 204.350 112.355 ;
        RECT 204.410 112.095 204.670 112.355 ;
        RECT 204.730 112.095 204.990 112.355 ;
        RECT 205.050 112.095 205.310 112.355 ;
        RECT 205.370 112.095 205.630 112.355 ;
        RECT 205.690 112.095 205.950 112.355 ;
        RECT 206.010 112.095 206.270 112.355 ;
        RECT 206.330 112.095 206.590 112.355 ;
        RECT 206.650 112.095 206.910 112.355 ;
        RECT 206.970 112.095 207.230 112.355 ;
        RECT 207.290 112.095 207.550 112.355 ;
        RECT 207.610 112.095 207.870 112.355 ;
        RECT 207.930 112.095 208.190 112.355 ;
        RECT 208.250 112.095 208.510 112.355 ;
        RECT 208.570 112.095 208.830 112.355 ;
        RECT 208.890 112.095 209.150 112.355 ;
        RECT 202.490 87.625 203.070 106.125 ;
        RECT 205.455 105.600 206.035 106.180 ;
        RECT 205.455 102.710 206.035 103.290 ;
        RECT 205.445 99.905 206.025 100.485 ;
        RECT 205.455 94.530 206.035 95.110 ;
        RECT 205.460 87.925 206.040 92.025 ;
        RECT 202.155 79.590 203.695 81.770 ;
        RECT 205.375 80.600 207.235 81.820 ;
        RECT 202.155 71.530 203.695 77.550 ;
      LAYER met2 ;
        RECT 201.125 110.645 209.250 117.060 ;
        RECT 201.125 108.790 207.300 110.645 ;
        RECT 201.125 70.950 203.830 108.790 ;
        RECT 205.310 81.885 207.300 108.790 ;
        RECT 205.310 80.785 207.305 81.885 ;
        RECT 205.315 80.520 207.305 80.785 ;
      LAYER via2 ;
        RECT 201.595 116.620 201.875 116.900 ;
        RECT 201.995 116.620 202.275 116.900 ;
        RECT 202.395 116.620 202.675 116.900 ;
        RECT 202.795 116.620 203.075 116.900 ;
        RECT 206.120 116.620 206.400 116.900 ;
        RECT 206.520 116.620 206.800 116.900 ;
        RECT 206.920 116.620 207.200 116.900 ;
        RECT 207.320 116.620 207.600 116.900 ;
        RECT 201.595 116.175 201.875 116.455 ;
        RECT 201.995 116.175 202.275 116.455 ;
        RECT 202.395 116.175 202.675 116.455 ;
        RECT 202.795 116.175 203.075 116.455 ;
        RECT 206.120 116.150 206.400 116.430 ;
        RECT 206.520 116.150 206.800 116.430 ;
        RECT 206.920 116.150 207.200 116.430 ;
        RECT 207.320 116.150 207.600 116.430 ;
      LAYER met3 ;
        RECT 201.125 116.050 209.250 117.060 ;
      LAYER via3 ;
        RECT 201.575 116.600 201.895 116.920 ;
        RECT 201.975 116.600 202.295 116.920 ;
        RECT 202.375 116.600 202.695 116.920 ;
        RECT 202.775 116.600 203.095 116.920 ;
        RECT 206.100 116.600 206.420 116.920 ;
        RECT 206.500 116.600 206.820 116.920 ;
        RECT 206.900 116.600 207.220 116.920 ;
        RECT 207.300 116.600 207.620 116.920 ;
        RECT 201.575 116.155 201.895 116.475 ;
        RECT 201.975 116.155 202.295 116.475 ;
        RECT 202.375 116.155 202.695 116.475 ;
        RECT 202.775 116.155 203.095 116.475 ;
        RECT 206.100 116.130 206.420 116.450 ;
        RECT 206.500 116.130 206.820 116.450 ;
        RECT 206.900 116.130 207.220 116.450 ;
        RECT 207.300 116.130 207.620 116.450 ;
      LAYER met4 ;
        RECT 201.565 0.000 203.165 211.800 ;
        RECT 206.090 0.000 207.690 211.800 ;
    END
  END vssa1
  OBS
      LAYER pwell ;
        RECT 202.720 71.690 203.460 77.720 ;
        RECT 227.000 71.690 227.740 77.720 ;
      LAYER li1 ;
        RECT 224.840 114.190 227.000 114.540 ;
        RECT 210.560 113.405 212.720 113.755 ;
        RECT 214.840 113.360 217.000 113.710 ;
        RECT 224.840 113.360 227.000 113.710 ;
        RECT 214.840 112.530 217.000 112.880 ;
        RECT 224.840 112.530 227.000 112.880 ;
        RECT 214.840 111.700 217.000 112.050 ;
        RECT 224.840 111.700 227.000 112.050 ;
        RECT 214.840 110.870 217.000 111.220 ;
        RECT 224.840 110.870 227.000 111.220 ;
        RECT 214.840 110.040 217.000 110.390 ;
        RECT 224.840 110.040 227.000 110.390 ;
        RECT 214.840 109.210 217.000 109.560 ;
        RECT 224.840 109.210 227.000 109.560 ;
        RECT 214.840 108.380 217.000 108.730 ;
        RECT 224.840 108.380 227.000 108.730 ;
        RECT 210.750 107.480 210.920 107.980 ;
        RECT 211.810 107.480 211.980 107.980 ;
        RECT 214.840 107.550 217.000 107.900 ;
        RECT 224.840 107.550 227.000 107.900 ;
        RECT 211.135 107.250 211.595 107.420 ;
        RECT 214.840 106.720 217.000 107.070 ;
        RECT 224.840 106.720 227.000 107.070 ;
        RECT 207.020 105.480 207.480 105.650 ;
        RECT 203.680 104.920 203.850 105.420 ;
        RECT 204.650 104.920 204.820 105.420 ;
        RECT 206.680 104.920 206.850 105.420 ;
        RECT 207.650 104.920 207.820 105.420 ;
        RECT 204.020 104.690 204.480 104.860 ;
        RECT 207.020 104.690 207.480 104.860 ;
        RECT 210.750 104.400 210.920 104.900 ;
        RECT 211.810 104.400 211.980 104.900 ;
        RECT 211.135 104.170 211.595 104.340 ;
        RECT 224.830 103.340 226.990 103.690 ;
        RECT 207.020 102.700 207.480 102.870 ;
        RECT 203.680 102.140 203.850 102.640 ;
        RECT 204.650 102.140 204.820 102.640 ;
        RECT 206.680 102.140 206.850 102.640 ;
        RECT 207.650 102.140 207.820 102.640 ;
        RECT 214.830 102.510 216.990 102.860 ;
        RECT 224.830 102.510 226.990 102.860 ;
        RECT 204.020 101.910 204.480 102.080 ;
        RECT 207.020 101.910 207.480 102.080 ;
        RECT 210.750 101.320 210.920 101.820 ;
        RECT 211.810 101.320 211.980 101.820 ;
        RECT 214.830 101.680 216.990 102.030 ;
        RECT 224.830 101.680 226.990 102.030 ;
        RECT 211.135 101.090 211.595 101.260 ;
        RECT 214.830 100.850 216.990 101.200 ;
        RECT 224.830 100.850 226.990 101.200 ;
        RECT 207.020 99.920 207.480 100.090 ;
        RECT 214.830 100.020 216.990 100.370 ;
        RECT 224.830 100.020 226.990 100.370 ;
        RECT 203.680 99.360 203.850 99.860 ;
        RECT 204.650 99.360 204.820 99.860 ;
        RECT 204.020 99.130 204.480 99.300 ;
        RECT 207.020 99.130 207.480 99.300 ;
        RECT 214.830 99.190 216.990 99.540 ;
        RECT 224.830 99.190 226.990 99.540 ;
        RECT 211.135 98.800 211.595 98.970 ;
        RECT 214.830 98.360 216.990 98.710 ;
        RECT 224.830 98.360 226.990 98.710 ;
        RECT 211.135 98.010 211.595 98.180 ;
        RECT 214.830 97.530 216.990 97.880 ;
        RECT 224.830 97.530 226.990 97.880 ;
        RECT 204.020 97.140 204.480 97.310 ;
        RECT 203.680 96.580 203.850 97.080 ;
        RECT 204.650 96.580 204.820 97.080 ;
        RECT 214.830 96.700 216.990 97.050 ;
        RECT 224.830 96.700 226.990 97.050 ;
        RECT 214.830 95.870 216.990 96.220 ;
        RECT 224.830 95.870 226.990 96.220 ;
        RECT 210.750 95.160 210.920 95.660 ;
        RECT 211.810 95.160 211.980 95.660 ;
        RECT 211.135 94.930 211.595 95.100 ;
        RECT 214.830 95.040 216.990 95.390 ;
        RECT 224.830 95.040 226.990 95.390 ;
        RECT 203.680 93.800 203.850 94.300 ;
        RECT 204.650 93.800 204.820 94.300 ;
        RECT 206.680 93.800 206.850 94.300 ;
        RECT 207.650 93.800 207.820 94.300 ;
        RECT 214.830 94.210 216.990 94.560 ;
        RECT 224.830 94.210 226.990 94.560 ;
        RECT 204.020 93.570 204.480 93.740 ;
        RECT 207.020 93.570 207.480 93.740 ;
        RECT 214.830 93.380 216.990 93.730 ;
        RECT 224.830 93.380 226.990 93.730 ;
        RECT 210.750 92.080 210.920 92.580 ;
        RECT 211.810 92.080 211.980 92.580 ;
        RECT 214.830 92.550 216.990 92.900 ;
        RECT 224.830 92.550 226.990 92.900 ;
        RECT 211.135 91.850 211.595 92.020 ;
        RECT 214.830 91.720 216.990 92.070 ;
        RECT 224.830 91.720 226.990 92.070 ;
        RECT 203.680 91.020 203.850 91.520 ;
        RECT 204.650 91.020 204.820 91.520 ;
        RECT 206.680 91.020 206.850 91.520 ;
        RECT 207.650 91.020 207.820 91.520 ;
        RECT 204.020 90.790 204.480 90.960 ;
        RECT 207.020 90.790 207.480 90.960 ;
        RECT 214.830 90.890 216.990 91.240 ;
        RECT 224.830 90.890 226.990 91.240 ;
        RECT 214.830 90.060 216.990 90.410 ;
        RECT 224.830 90.060 226.990 90.410 ;
        RECT 210.750 89.000 210.920 89.500 ;
        RECT 211.810 89.000 211.980 89.500 ;
        RECT 214.830 89.230 216.990 89.580 ;
        RECT 224.830 89.230 226.990 89.580 ;
        RECT 204.020 88.800 204.480 88.970 ;
        RECT 211.135 88.770 211.595 88.940 ;
        RECT 203.680 88.240 203.850 88.740 ;
        RECT 204.650 88.240 204.820 88.740 ;
        RECT 206.680 88.240 206.850 88.740 ;
        RECT 207.650 88.240 207.820 88.740 ;
        RECT 214.830 88.400 216.990 88.750 ;
        RECT 224.830 88.400 226.990 88.750 ;
        RECT 204.020 88.010 204.480 88.180 ;
        RECT 207.020 88.010 207.480 88.180 ;
        RECT 214.830 87.570 216.990 87.920 ;
        RECT 224.830 87.570 226.990 87.920 ;
        RECT 214.830 86.740 216.990 87.090 ;
        RECT 224.830 86.740 226.990 87.090 ;
        RECT 211.135 86.480 211.595 86.650 ;
        RECT 210.750 85.920 210.920 86.420 ;
        RECT 211.810 85.920 211.980 86.420 ;
        RECT 214.830 85.910 216.990 86.260 ;
        RECT 224.830 85.910 226.990 86.260 ;
        RECT 211.135 85.690 211.595 85.860 ;
        RECT 214.830 85.080 216.990 85.430 ;
        RECT 224.830 85.080 226.990 85.430 ;
        RECT 214.830 84.250 216.990 84.600 ;
        RECT 224.830 84.250 226.990 84.600 ;
        RECT 203.545 83.195 205.705 83.545 ;
        RECT 210.545 83.195 212.705 83.545 ;
        RECT 214.830 83.420 216.990 83.770 ;
        RECT 224.830 83.420 226.990 83.770 ;
        RECT 203.545 82.365 205.705 82.715 ;
        RECT 212.830 80.180 214.990 80.530 ;
        RECT 202.850 71.860 203.330 77.550 ;
        RECT 208.895 76.360 209.355 76.530 ;
        RECT 212.245 76.360 212.705 76.530 ;
        RECT 217.755 76.360 218.215 76.530 ;
        RECT 221.105 76.360 221.565 76.530 ;
        RECT 205.060 75.790 205.230 76.290 ;
        RECT 206.030 75.790 206.200 76.290 ;
        RECT 208.510 75.800 208.680 76.300 ;
        RECT 209.570 75.800 209.740 76.300 ;
        RECT 211.860 75.800 212.030 76.300 ;
        RECT 212.920 75.800 213.090 76.300 ;
        RECT 217.370 75.800 217.540 76.300 ;
        RECT 218.430 75.800 218.600 76.300 ;
        RECT 220.720 75.800 220.890 76.300 ;
        RECT 221.780 75.800 221.950 76.300 ;
        RECT 224.260 75.790 224.430 76.290 ;
        RECT 225.230 75.790 225.400 76.290 ;
        RECT 205.400 75.560 205.860 75.730 ;
        RECT 208.895 75.570 209.355 75.740 ;
        RECT 221.105 75.570 221.565 75.740 ;
        RECT 224.600 75.560 225.060 75.730 ;
        RECT 205.390 73.320 205.850 73.490 ;
        RECT 208.905 73.310 209.365 73.480 ;
        RECT 221.095 73.310 221.555 73.480 ;
        RECT 224.610 73.320 225.070 73.490 ;
        RECT 208.520 72.750 208.690 73.250 ;
        RECT 209.580 72.750 209.750 73.250 ;
        RECT 211.860 72.720 212.030 73.220 ;
        RECT 212.920 72.720 213.090 73.220 ;
        RECT 217.370 72.720 217.540 73.220 ;
        RECT 218.430 72.720 218.600 73.220 ;
        RECT 220.710 72.750 220.880 73.250 ;
        RECT 221.770 72.750 221.940 73.250 ;
        RECT 208.905 72.520 209.365 72.690 ;
        RECT 212.245 72.490 212.705 72.660 ;
        RECT 217.755 72.490 218.215 72.660 ;
        RECT 221.095 72.520 221.555 72.690 ;
        RECT 227.130 71.860 227.610 77.550 ;
        RECT 213.880 65.350 214.210 65.520 ;
        RECT 206.720 64.870 207.760 65.040 ;
        RECT 209.910 64.870 210.950 65.040 ;
        RECT 216.250 64.905 216.580 65.075 ;
        RECT 219.510 64.870 220.550 65.040 ;
        RECT 222.700 64.870 223.740 65.040 ;
      LAYER mcon ;
        RECT 224.930 114.280 225.100 114.450 ;
        RECT 225.290 114.280 225.460 114.450 ;
        RECT 225.650 114.280 225.820 114.450 ;
        RECT 226.010 114.280 226.180 114.450 ;
        RECT 226.370 114.280 226.540 114.450 ;
        RECT 226.730 114.280 226.900 114.450 ;
        RECT 210.650 113.495 210.820 113.665 ;
        RECT 211.010 113.495 211.180 113.665 ;
        RECT 211.370 113.495 211.540 113.665 ;
        RECT 211.730 113.495 211.900 113.665 ;
        RECT 212.090 113.495 212.260 113.665 ;
        RECT 212.450 113.495 212.620 113.665 ;
        RECT 214.935 113.450 215.105 113.620 ;
        RECT 215.295 113.450 215.465 113.620 ;
        RECT 215.655 113.450 215.825 113.620 ;
        RECT 216.015 113.450 216.185 113.620 ;
        RECT 216.375 113.450 216.545 113.620 ;
        RECT 216.735 113.450 216.905 113.620 ;
        RECT 224.930 113.450 225.100 113.620 ;
        RECT 225.290 113.450 225.460 113.620 ;
        RECT 225.650 113.450 225.820 113.620 ;
        RECT 226.010 113.450 226.180 113.620 ;
        RECT 226.370 113.450 226.540 113.620 ;
        RECT 226.730 113.450 226.900 113.620 ;
        RECT 214.935 112.620 215.105 112.790 ;
        RECT 215.295 112.620 215.465 112.790 ;
        RECT 215.655 112.620 215.825 112.790 ;
        RECT 216.015 112.620 216.185 112.790 ;
        RECT 216.375 112.620 216.545 112.790 ;
        RECT 216.735 112.620 216.905 112.790 ;
        RECT 224.930 112.620 225.100 112.790 ;
        RECT 225.290 112.620 225.460 112.790 ;
        RECT 225.650 112.620 225.820 112.790 ;
        RECT 226.010 112.620 226.180 112.790 ;
        RECT 226.370 112.620 226.540 112.790 ;
        RECT 226.730 112.620 226.900 112.790 ;
        RECT 214.935 111.790 215.105 111.960 ;
        RECT 215.295 111.790 215.465 111.960 ;
        RECT 215.655 111.790 215.825 111.960 ;
        RECT 216.015 111.790 216.185 111.960 ;
        RECT 216.375 111.790 216.545 111.960 ;
        RECT 216.735 111.790 216.905 111.960 ;
        RECT 224.930 111.790 225.100 111.960 ;
        RECT 225.290 111.790 225.460 111.960 ;
        RECT 225.650 111.790 225.820 111.960 ;
        RECT 226.010 111.790 226.180 111.960 ;
        RECT 226.370 111.790 226.540 111.960 ;
        RECT 226.730 111.790 226.900 111.960 ;
        RECT 214.935 110.960 215.105 111.130 ;
        RECT 215.295 110.960 215.465 111.130 ;
        RECT 215.655 110.960 215.825 111.130 ;
        RECT 216.015 110.960 216.185 111.130 ;
        RECT 216.375 110.960 216.545 111.130 ;
        RECT 216.735 110.960 216.905 111.130 ;
        RECT 224.930 110.960 225.100 111.130 ;
        RECT 225.290 110.960 225.460 111.130 ;
        RECT 225.650 110.960 225.820 111.130 ;
        RECT 226.010 110.960 226.180 111.130 ;
        RECT 226.370 110.960 226.540 111.130 ;
        RECT 226.730 110.960 226.900 111.130 ;
        RECT 214.935 110.130 215.105 110.300 ;
        RECT 215.295 110.130 215.465 110.300 ;
        RECT 215.655 110.130 215.825 110.300 ;
        RECT 216.015 110.130 216.185 110.300 ;
        RECT 216.375 110.130 216.545 110.300 ;
        RECT 216.735 110.130 216.905 110.300 ;
        RECT 224.930 110.130 225.100 110.300 ;
        RECT 225.290 110.130 225.460 110.300 ;
        RECT 225.650 110.130 225.820 110.300 ;
        RECT 226.010 110.130 226.180 110.300 ;
        RECT 226.370 110.130 226.540 110.300 ;
        RECT 226.730 110.130 226.900 110.300 ;
        RECT 214.935 109.300 215.105 109.470 ;
        RECT 215.295 109.300 215.465 109.470 ;
        RECT 215.655 109.300 215.825 109.470 ;
        RECT 216.015 109.300 216.185 109.470 ;
        RECT 216.375 109.300 216.545 109.470 ;
        RECT 216.735 109.300 216.905 109.470 ;
        RECT 224.930 109.300 225.100 109.470 ;
        RECT 225.290 109.300 225.460 109.470 ;
        RECT 225.650 109.300 225.820 109.470 ;
        RECT 226.010 109.300 226.180 109.470 ;
        RECT 226.370 109.300 226.540 109.470 ;
        RECT 226.730 109.300 226.900 109.470 ;
        RECT 214.935 108.470 215.105 108.640 ;
        RECT 215.295 108.470 215.465 108.640 ;
        RECT 215.655 108.470 215.825 108.640 ;
        RECT 216.015 108.470 216.185 108.640 ;
        RECT 216.375 108.470 216.545 108.640 ;
        RECT 216.735 108.470 216.905 108.640 ;
        RECT 224.930 108.470 225.100 108.640 ;
        RECT 225.290 108.470 225.460 108.640 ;
        RECT 225.650 108.470 225.820 108.640 ;
        RECT 226.010 108.470 226.180 108.640 ;
        RECT 226.370 108.470 226.540 108.640 ;
        RECT 226.730 108.470 226.900 108.640 ;
        RECT 210.750 107.645 210.920 107.815 ;
        RECT 211.810 107.645 211.980 107.815 ;
        RECT 214.935 107.640 215.105 107.810 ;
        RECT 215.295 107.640 215.465 107.810 ;
        RECT 215.655 107.640 215.825 107.810 ;
        RECT 216.015 107.640 216.185 107.810 ;
        RECT 216.375 107.640 216.545 107.810 ;
        RECT 216.735 107.640 216.905 107.810 ;
        RECT 224.930 107.640 225.100 107.810 ;
        RECT 225.290 107.640 225.460 107.810 ;
        RECT 225.650 107.640 225.820 107.810 ;
        RECT 226.010 107.640 226.180 107.810 ;
        RECT 226.370 107.640 226.540 107.810 ;
        RECT 226.730 107.640 226.900 107.810 ;
        RECT 211.280 107.250 211.450 107.420 ;
        RECT 214.935 106.810 215.105 106.980 ;
        RECT 215.295 106.810 215.465 106.980 ;
        RECT 215.655 106.810 215.825 106.980 ;
        RECT 216.015 106.810 216.185 106.980 ;
        RECT 216.375 106.810 216.545 106.980 ;
        RECT 216.735 106.810 216.905 106.980 ;
        RECT 224.930 106.810 225.100 106.980 ;
        RECT 225.290 106.810 225.460 106.980 ;
        RECT 225.650 106.810 225.820 106.980 ;
        RECT 226.010 106.810 226.180 106.980 ;
        RECT 226.370 106.810 226.540 106.980 ;
        RECT 226.730 106.810 226.900 106.980 ;
        RECT 207.165 105.480 207.335 105.650 ;
        RECT 203.680 105.085 203.850 105.255 ;
        RECT 204.650 105.085 204.820 105.255 ;
        RECT 206.680 105.085 206.850 105.255 ;
        RECT 207.650 105.085 207.820 105.255 ;
        RECT 204.165 104.690 204.335 104.860 ;
        RECT 207.165 104.690 207.335 104.860 ;
        RECT 210.750 104.565 210.920 104.735 ;
        RECT 211.810 104.565 211.980 104.735 ;
        RECT 211.280 104.170 211.450 104.340 ;
        RECT 224.920 103.430 225.090 103.600 ;
        RECT 225.280 103.430 225.450 103.600 ;
        RECT 225.640 103.430 225.810 103.600 ;
        RECT 226.000 103.430 226.170 103.600 ;
        RECT 226.360 103.430 226.530 103.600 ;
        RECT 226.720 103.430 226.890 103.600 ;
        RECT 207.165 102.700 207.335 102.870 ;
        RECT 203.680 102.305 203.850 102.475 ;
        RECT 204.650 102.305 204.820 102.475 ;
        RECT 206.680 102.305 206.850 102.475 ;
        RECT 214.925 102.600 215.095 102.770 ;
        RECT 215.285 102.600 215.455 102.770 ;
        RECT 215.645 102.600 215.815 102.770 ;
        RECT 216.005 102.600 216.175 102.770 ;
        RECT 216.365 102.600 216.535 102.770 ;
        RECT 216.725 102.600 216.895 102.770 ;
        RECT 224.920 102.600 225.090 102.770 ;
        RECT 225.280 102.600 225.450 102.770 ;
        RECT 225.640 102.600 225.810 102.770 ;
        RECT 226.000 102.600 226.170 102.770 ;
        RECT 226.360 102.600 226.530 102.770 ;
        RECT 226.720 102.600 226.890 102.770 ;
        RECT 207.650 102.305 207.820 102.475 ;
        RECT 204.165 101.910 204.335 102.080 ;
        RECT 207.165 101.910 207.335 102.080 ;
        RECT 210.750 101.485 210.920 101.655 ;
        RECT 214.925 101.770 215.095 101.940 ;
        RECT 215.285 101.770 215.455 101.940 ;
        RECT 215.645 101.770 215.815 101.940 ;
        RECT 216.005 101.770 216.175 101.940 ;
        RECT 216.365 101.770 216.535 101.940 ;
        RECT 216.725 101.770 216.895 101.940 ;
        RECT 224.920 101.770 225.090 101.940 ;
        RECT 225.280 101.770 225.450 101.940 ;
        RECT 225.640 101.770 225.810 101.940 ;
        RECT 226.000 101.770 226.170 101.940 ;
        RECT 226.360 101.770 226.530 101.940 ;
        RECT 226.720 101.770 226.890 101.940 ;
        RECT 211.810 101.485 211.980 101.655 ;
        RECT 211.280 101.090 211.450 101.260 ;
        RECT 214.925 100.940 215.095 101.110 ;
        RECT 215.285 100.940 215.455 101.110 ;
        RECT 215.645 100.940 215.815 101.110 ;
        RECT 216.005 100.940 216.175 101.110 ;
        RECT 216.365 100.940 216.535 101.110 ;
        RECT 216.725 100.940 216.895 101.110 ;
        RECT 224.920 100.940 225.090 101.110 ;
        RECT 225.280 100.940 225.450 101.110 ;
        RECT 225.640 100.940 225.810 101.110 ;
        RECT 226.000 100.940 226.170 101.110 ;
        RECT 226.360 100.940 226.530 101.110 ;
        RECT 226.720 100.940 226.890 101.110 ;
        RECT 214.925 100.110 215.095 100.280 ;
        RECT 215.285 100.110 215.455 100.280 ;
        RECT 215.645 100.110 215.815 100.280 ;
        RECT 216.005 100.110 216.175 100.280 ;
        RECT 216.365 100.110 216.535 100.280 ;
        RECT 216.725 100.110 216.895 100.280 ;
        RECT 207.165 99.920 207.335 100.090 ;
        RECT 224.920 100.110 225.090 100.280 ;
        RECT 225.280 100.110 225.450 100.280 ;
        RECT 225.640 100.110 225.810 100.280 ;
        RECT 226.000 100.110 226.170 100.280 ;
        RECT 226.360 100.110 226.530 100.280 ;
        RECT 226.720 100.110 226.890 100.280 ;
        RECT 203.680 99.525 203.850 99.695 ;
        RECT 204.650 99.525 204.820 99.695 ;
        RECT 204.165 99.130 204.335 99.300 ;
        RECT 207.165 99.130 207.335 99.300 ;
        RECT 214.925 99.280 215.095 99.450 ;
        RECT 215.285 99.280 215.455 99.450 ;
        RECT 215.645 99.280 215.815 99.450 ;
        RECT 216.005 99.280 216.175 99.450 ;
        RECT 216.365 99.280 216.535 99.450 ;
        RECT 216.725 99.280 216.895 99.450 ;
        RECT 224.920 99.280 225.090 99.450 ;
        RECT 225.280 99.280 225.450 99.450 ;
        RECT 225.640 99.280 225.810 99.450 ;
        RECT 226.000 99.280 226.170 99.450 ;
        RECT 226.360 99.280 226.530 99.450 ;
        RECT 226.720 99.280 226.890 99.450 ;
        RECT 211.280 98.800 211.450 98.970 ;
        RECT 214.925 98.450 215.095 98.620 ;
        RECT 215.285 98.450 215.455 98.620 ;
        RECT 215.645 98.450 215.815 98.620 ;
        RECT 216.005 98.450 216.175 98.620 ;
        RECT 216.365 98.450 216.535 98.620 ;
        RECT 216.725 98.450 216.895 98.620 ;
        RECT 224.920 98.450 225.090 98.620 ;
        RECT 225.280 98.450 225.450 98.620 ;
        RECT 225.640 98.450 225.810 98.620 ;
        RECT 226.000 98.450 226.170 98.620 ;
        RECT 226.360 98.450 226.530 98.620 ;
        RECT 226.720 98.450 226.890 98.620 ;
        RECT 211.280 98.010 211.450 98.180 ;
        RECT 214.925 97.620 215.095 97.790 ;
        RECT 215.285 97.620 215.455 97.790 ;
        RECT 215.645 97.620 215.815 97.790 ;
        RECT 216.005 97.620 216.175 97.790 ;
        RECT 216.365 97.620 216.535 97.790 ;
        RECT 216.725 97.620 216.895 97.790 ;
        RECT 224.920 97.620 225.090 97.790 ;
        RECT 225.280 97.620 225.450 97.790 ;
        RECT 225.640 97.620 225.810 97.790 ;
        RECT 226.000 97.620 226.170 97.790 ;
        RECT 226.360 97.620 226.530 97.790 ;
        RECT 226.720 97.620 226.890 97.790 ;
        RECT 204.165 97.140 204.335 97.310 ;
        RECT 203.680 96.745 203.850 96.915 ;
        RECT 204.650 96.745 204.820 96.915 ;
        RECT 214.925 96.790 215.095 96.960 ;
        RECT 215.285 96.790 215.455 96.960 ;
        RECT 215.645 96.790 215.815 96.960 ;
        RECT 216.005 96.790 216.175 96.960 ;
        RECT 216.365 96.790 216.535 96.960 ;
        RECT 216.725 96.790 216.895 96.960 ;
        RECT 224.920 96.790 225.090 96.960 ;
        RECT 225.280 96.790 225.450 96.960 ;
        RECT 225.640 96.790 225.810 96.960 ;
        RECT 226.000 96.790 226.170 96.960 ;
        RECT 226.360 96.790 226.530 96.960 ;
        RECT 226.720 96.790 226.890 96.960 ;
        RECT 214.925 95.960 215.095 96.130 ;
        RECT 215.285 95.960 215.455 96.130 ;
        RECT 215.645 95.960 215.815 96.130 ;
        RECT 216.005 95.960 216.175 96.130 ;
        RECT 216.365 95.960 216.535 96.130 ;
        RECT 216.725 95.960 216.895 96.130 ;
        RECT 224.920 95.960 225.090 96.130 ;
        RECT 225.280 95.960 225.450 96.130 ;
        RECT 225.640 95.960 225.810 96.130 ;
        RECT 226.000 95.960 226.170 96.130 ;
        RECT 226.360 95.960 226.530 96.130 ;
        RECT 226.720 95.960 226.890 96.130 ;
        RECT 210.750 95.325 210.920 95.495 ;
        RECT 211.810 95.325 211.980 95.495 ;
        RECT 214.925 95.130 215.095 95.300 ;
        RECT 215.285 95.130 215.455 95.300 ;
        RECT 215.645 95.130 215.815 95.300 ;
        RECT 216.005 95.130 216.175 95.300 ;
        RECT 216.365 95.130 216.535 95.300 ;
        RECT 216.725 95.130 216.895 95.300 ;
        RECT 211.280 94.930 211.450 95.100 ;
        RECT 224.920 95.130 225.090 95.300 ;
        RECT 225.280 95.130 225.450 95.300 ;
        RECT 225.640 95.130 225.810 95.300 ;
        RECT 226.000 95.130 226.170 95.300 ;
        RECT 226.360 95.130 226.530 95.300 ;
        RECT 226.720 95.130 226.890 95.300 ;
        RECT 214.925 94.300 215.095 94.470 ;
        RECT 215.285 94.300 215.455 94.470 ;
        RECT 215.645 94.300 215.815 94.470 ;
        RECT 216.005 94.300 216.175 94.470 ;
        RECT 216.365 94.300 216.535 94.470 ;
        RECT 216.725 94.300 216.895 94.470 ;
        RECT 203.680 93.965 203.850 94.135 ;
        RECT 204.650 93.965 204.820 94.135 ;
        RECT 206.680 93.965 206.850 94.135 ;
        RECT 224.920 94.300 225.090 94.470 ;
        RECT 225.280 94.300 225.450 94.470 ;
        RECT 225.640 94.300 225.810 94.470 ;
        RECT 226.000 94.300 226.170 94.470 ;
        RECT 226.360 94.300 226.530 94.470 ;
        RECT 226.720 94.300 226.890 94.470 ;
        RECT 207.650 93.965 207.820 94.135 ;
        RECT 204.165 93.570 204.335 93.740 ;
        RECT 207.165 93.570 207.335 93.740 ;
        RECT 214.925 93.470 215.095 93.640 ;
        RECT 215.285 93.470 215.455 93.640 ;
        RECT 215.645 93.470 215.815 93.640 ;
        RECT 216.005 93.470 216.175 93.640 ;
        RECT 216.365 93.470 216.535 93.640 ;
        RECT 216.725 93.470 216.895 93.640 ;
        RECT 224.920 93.470 225.090 93.640 ;
        RECT 225.280 93.470 225.450 93.640 ;
        RECT 225.640 93.470 225.810 93.640 ;
        RECT 226.000 93.470 226.170 93.640 ;
        RECT 226.360 93.470 226.530 93.640 ;
        RECT 226.720 93.470 226.890 93.640 ;
        RECT 214.925 92.640 215.095 92.810 ;
        RECT 215.285 92.640 215.455 92.810 ;
        RECT 215.645 92.640 215.815 92.810 ;
        RECT 216.005 92.640 216.175 92.810 ;
        RECT 216.365 92.640 216.535 92.810 ;
        RECT 216.725 92.640 216.895 92.810 ;
        RECT 210.750 92.245 210.920 92.415 ;
        RECT 224.920 92.640 225.090 92.810 ;
        RECT 225.280 92.640 225.450 92.810 ;
        RECT 225.640 92.640 225.810 92.810 ;
        RECT 226.000 92.640 226.170 92.810 ;
        RECT 226.360 92.640 226.530 92.810 ;
        RECT 226.720 92.640 226.890 92.810 ;
        RECT 211.810 92.245 211.980 92.415 ;
        RECT 211.280 91.850 211.450 92.020 ;
        RECT 214.925 91.810 215.095 91.980 ;
        RECT 215.285 91.810 215.455 91.980 ;
        RECT 215.645 91.810 215.815 91.980 ;
        RECT 216.005 91.810 216.175 91.980 ;
        RECT 216.365 91.810 216.535 91.980 ;
        RECT 216.725 91.810 216.895 91.980 ;
        RECT 224.920 91.810 225.090 91.980 ;
        RECT 225.280 91.810 225.450 91.980 ;
        RECT 225.640 91.810 225.810 91.980 ;
        RECT 226.000 91.810 226.170 91.980 ;
        RECT 226.360 91.810 226.530 91.980 ;
        RECT 226.720 91.810 226.890 91.980 ;
        RECT 203.680 91.185 203.850 91.355 ;
        RECT 204.650 91.185 204.820 91.355 ;
        RECT 206.680 91.185 206.850 91.355 ;
        RECT 207.650 91.185 207.820 91.355 ;
        RECT 214.925 90.980 215.095 91.150 ;
        RECT 215.285 90.980 215.455 91.150 ;
        RECT 215.645 90.980 215.815 91.150 ;
        RECT 216.005 90.980 216.175 91.150 ;
        RECT 216.365 90.980 216.535 91.150 ;
        RECT 216.725 90.980 216.895 91.150 ;
        RECT 204.165 90.790 204.335 90.960 ;
        RECT 207.165 90.790 207.335 90.960 ;
        RECT 224.920 90.980 225.090 91.150 ;
        RECT 225.280 90.980 225.450 91.150 ;
        RECT 225.640 90.980 225.810 91.150 ;
        RECT 226.000 90.980 226.170 91.150 ;
        RECT 226.360 90.980 226.530 91.150 ;
        RECT 226.720 90.980 226.890 91.150 ;
        RECT 214.925 90.150 215.095 90.320 ;
        RECT 215.285 90.150 215.455 90.320 ;
        RECT 215.645 90.150 215.815 90.320 ;
        RECT 216.005 90.150 216.175 90.320 ;
        RECT 216.365 90.150 216.535 90.320 ;
        RECT 216.725 90.150 216.895 90.320 ;
        RECT 224.920 90.150 225.090 90.320 ;
        RECT 225.280 90.150 225.450 90.320 ;
        RECT 225.640 90.150 225.810 90.320 ;
        RECT 226.000 90.150 226.170 90.320 ;
        RECT 226.360 90.150 226.530 90.320 ;
        RECT 226.720 90.150 226.890 90.320 ;
        RECT 210.750 89.165 210.920 89.335 ;
        RECT 211.810 89.165 211.980 89.335 ;
        RECT 214.925 89.320 215.095 89.490 ;
        RECT 215.285 89.320 215.455 89.490 ;
        RECT 215.645 89.320 215.815 89.490 ;
        RECT 216.005 89.320 216.175 89.490 ;
        RECT 216.365 89.320 216.535 89.490 ;
        RECT 216.725 89.320 216.895 89.490 ;
        RECT 224.920 89.320 225.090 89.490 ;
        RECT 225.280 89.320 225.450 89.490 ;
        RECT 225.640 89.320 225.810 89.490 ;
        RECT 226.000 89.320 226.170 89.490 ;
        RECT 226.360 89.320 226.530 89.490 ;
        RECT 226.720 89.320 226.890 89.490 ;
        RECT 204.165 88.800 204.335 88.970 ;
        RECT 211.280 88.770 211.450 88.940 ;
        RECT 203.680 88.405 203.850 88.575 ;
        RECT 204.650 88.405 204.820 88.575 ;
        RECT 206.680 88.405 206.850 88.575 ;
        RECT 207.650 88.405 207.820 88.575 ;
        RECT 214.925 88.490 215.095 88.660 ;
        RECT 215.285 88.490 215.455 88.660 ;
        RECT 215.645 88.490 215.815 88.660 ;
        RECT 216.005 88.490 216.175 88.660 ;
        RECT 216.365 88.490 216.535 88.660 ;
        RECT 216.725 88.490 216.895 88.660 ;
        RECT 224.920 88.490 225.090 88.660 ;
        RECT 225.280 88.490 225.450 88.660 ;
        RECT 225.640 88.490 225.810 88.660 ;
        RECT 226.000 88.490 226.170 88.660 ;
        RECT 226.360 88.490 226.530 88.660 ;
        RECT 226.720 88.490 226.890 88.660 ;
        RECT 204.165 88.010 204.335 88.180 ;
        RECT 207.165 88.010 207.335 88.180 ;
        RECT 214.925 87.660 215.095 87.830 ;
        RECT 215.285 87.660 215.455 87.830 ;
        RECT 215.645 87.660 215.815 87.830 ;
        RECT 216.005 87.660 216.175 87.830 ;
        RECT 216.365 87.660 216.535 87.830 ;
        RECT 216.725 87.660 216.895 87.830 ;
        RECT 224.920 87.660 225.090 87.830 ;
        RECT 225.280 87.660 225.450 87.830 ;
        RECT 225.640 87.660 225.810 87.830 ;
        RECT 226.000 87.660 226.170 87.830 ;
        RECT 226.360 87.660 226.530 87.830 ;
        RECT 226.720 87.660 226.890 87.830 ;
        RECT 214.925 86.830 215.095 87.000 ;
        RECT 215.285 86.830 215.455 87.000 ;
        RECT 215.645 86.830 215.815 87.000 ;
        RECT 216.005 86.830 216.175 87.000 ;
        RECT 216.365 86.830 216.535 87.000 ;
        RECT 216.725 86.830 216.895 87.000 ;
        RECT 224.920 86.830 225.090 87.000 ;
        RECT 225.280 86.830 225.450 87.000 ;
        RECT 225.640 86.830 225.810 87.000 ;
        RECT 226.000 86.830 226.170 87.000 ;
        RECT 226.360 86.830 226.530 87.000 ;
        RECT 226.720 86.830 226.890 87.000 ;
        RECT 211.280 86.480 211.450 86.650 ;
        RECT 210.750 86.085 210.920 86.255 ;
        RECT 211.810 86.085 211.980 86.255 ;
        RECT 214.925 86.000 215.095 86.170 ;
        RECT 215.285 86.000 215.455 86.170 ;
        RECT 215.645 86.000 215.815 86.170 ;
        RECT 216.005 86.000 216.175 86.170 ;
        RECT 216.365 86.000 216.535 86.170 ;
        RECT 216.725 86.000 216.895 86.170 ;
        RECT 224.920 86.000 225.090 86.170 ;
        RECT 225.280 86.000 225.450 86.170 ;
        RECT 225.640 86.000 225.810 86.170 ;
        RECT 226.000 86.000 226.170 86.170 ;
        RECT 226.360 86.000 226.530 86.170 ;
        RECT 226.720 86.000 226.890 86.170 ;
        RECT 211.280 85.690 211.450 85.860 ;
        RECT 214.925 85.170 215.095 85.340 ;
        RECT 215.285 85.170 215.455 85.340 ;
        RECT 215.645 85.170 215.815 85.340 ;
        RECT 216.005 85.170 216.175 85.340 ;
        RECT 216.365 85.170 216.535 85.340 ;
        RECT 216.725 85.170 216.895 85.340 ;
        RECT 224.920 85.170 225.090 85.340 ;
        RECT 225.280 85.170 225.450 85.340 ;
        RECT 225.640 85.170 225.810 85.340 ;
        RECT 226.000 85.170 226.170 85.340 ;
        RECT 226.360 85.170 226.530 85.340 ;
        RECT 226.720 85.170 226.890 85.340 ;
        RECT 214.925 84.340 215.095 84.510 ;
        RECT 215.285 84.340 215.455 84.510 ;
        RECT 215.645 84.340 215.815 84.510 ;
        RECT 216.005 84.340 216.175 84.510 ;
        RECT 216.365 84.340 216.535 84.510 ;
        RECT 216.725 84.340 216.895 84.510 ;
        RECT 224.920 84.340 225.090 84.510 ;
        RECT 225.280 84.340 225.450 84.510 ;
        RECT 225.640 84.340 225.810 84.510 ;
        RECT 226.000 84.340 226.170 84.510 ;
        RECT 226.360 84.340 226.530 84.510 ;
        RECT 226.720 84.340 226.890 84.510 ;
        RECT 203.640 83.285 203.810 83.455 ;
        RECT 204.000 83.285 204.170 83.455 ;
        RECT 204.360 83.285 204.530 83.455 ;
        RECT 204.720 83.285 204.890 83.455 ;
        RECT 205.080 83.285 205.250 83.455 ;
        RECT 205.440 83.285 205.610 83.455 ;
        RECT 210.635 83.285 210.805 83.455 ;
        RECT 210.995 83.285 211.165 83.455 ;
        RECT 211.355 83.285 211.525 83.455 ;
        RECT 211.715 83.285 211.885 83.455 ;
        RECT 212.075 83.285 212.245 83.455 ;
        RECT 212.435 83.285 212.605 83.455 ;
        RECT 214.925 83.510 215.095 83.680 ;
        RECT 215.285 83.510 215.455 83.680 ;
        RECT 215.645 83.510 215.815 83.680 ;
        RECT 216.005 83.510 216.175 83.680 ;
        RECT 216.365 83.510 216.535 83.680 ;
        RECT 216.725 83.510 216.895 83.680 ;
        RECT 224.920 83.510 225.090 83.680 ;
        RECT 225.280 83.510 225.450 83.680 ;
        RECT 225.640 83.510 225.810 83.680 ;
        RECT 226.000 83.510 226.170 83.680 ;
        RECT 226.360 83.510 226.530 83.680 ;
        RECT 226.720 83.510 226.890 83.680 ;
        RECT 203.640 82.455 203.810 82.625 ;
        RECT 204.000 82.455 204.170 82.625 ;
        RECT 204.360 82.455 204.530 82.625 ;
        RECT 204.720 82.455 204.890 82.625 ;
        RECT 205.080 82.455 205.250 82.625 ;
        RECT 205.440 82.455 205.610 82.625 ;
        RECT 212.925 80.270 213.095 80.440 ;
        RECT 213.285 80.270 213.455 80.440 ;
        RECT 213.645 80.270 213.815 80.440 ;
        RECT 214.005 80.270 214.175 80.440 ;
        RECT 214.365 80.270 214.535 80.440 ;
        RECT 214.725 80.270 214.895 80.440 ;
        RECT 209.040 76.360 209.210 76.530 ;
        RECT 212.390 76.360 212.560 76.530 ;
        RECT 217.900 76.360 218.070 76.530 ;
        RECT 221.250 76.360 221.420 76.530 ;
        RECT 205.060 75.955 205.230 76.125 ;
        RECT 206.030 75.955 206.200 76.125 ;
        RECT 208.510 75.965 208.680 76.135 ;
        RECT 209.570 75.965 209.740 76.135 ;
        RECT 211.860 75.965 212.030 76.135 ;
        RECT 212.920 75.965 213.090 76.135 ;
        RECT 217.370 75.965 217.540 76.135 ;
        RECT 218.430 75.965 218.600 76.135 ;
        RECT 220.720 75.965 220.890 76.135 ;
        RECT 221.780 75.965 221.950 76.135 ;
        RECT 224.260 75.955 224.430 76.125 ;
        RECT 225.230 75.955 225.400 76.125 ;
        RECT 205.545 75.560 205.715 75.730 ;
        RECT 209.040 75.570 209.210 75.740 ;
        RECT 221.250 75.570 221.420 75.740 ;
        RECT 224.745 75.560 224.915 75.730 ;
        RECT 205.535 73.320 205.705 73.490 ;
        RECT 209.050 73.310 209.220 73.480 ;
        RECT 221.240 73.310 221.410 73.480 ;
        RECT 224.755 73.320 224.925 73.490 ;
        RECT 208.520 72.915 208.690 73.085 ;
        RECT 209.580 72.915 209.750 73.085 ;
        RECT 211.860 72.885 212.030 73.055 ;
        RECT 212.920 72.885 213.090 73.055 ;
        RECT 217.370 72.885 217.540 73.055 ;
        RECT 218.430 72.885 218.600 73.055 ;
        RECT 220.710 72.915 220.880 73.085 ;
        RECT 221.770 72.915 221.940 73.085 ;
        RECT 209.050 72.520 209.220 72.690 ;
        RECT 212.390 72.490 212.560 72.660 ;
        RECT 217.900 72.490 218.070 72.660 ;
        RECT 221.240 72.520 221.410 72.690 ;
        RECT 213.960 65.350 214.130 65.520 ;
        RECT 206.975 64.870 207.145 65.040 ;
        RECT 207.335 64.870 207.505 65.040 ;
        RECT 210.165 64.870 210.335 65.040 ;
        RECT 210.525 64.870 210.695 65.040 ;
        RECT 216.330 64.905 216.500 65.075 ;
        RECT 219.765 64.870 219.935 65.040 ;
        RECT 220.125 64.870 220.295 65.040 ;
        RECT 222.955 64.870 223.125 65.040 ;
        RECT 223.315 64.870 223.485 65.040 ;
      LAYER met1 ;
        RECT 210.585 113.680 212.690 113.705 ;
        RECT 213.895 113.680 214.220 113.880 ;
        RECT 210.585 113.465 214.220 113.680 ;
        RECT 210.585 113.455 212.690 113.465 ;
        RECT 213.895 112.775 214.220 113.465 ;
        RECT 214.840 112.530 217.000 113.710 ;
        RECT 224.840 113.360 227.000 114.540 ;
        RECT 214.840 110.870 217.000 112.050 ;
        RECT 224.840 111.700 227.000 112.880 ;
        RECT 207.180 109.440 213.810 109.625 ;
        RECT 207.180 105.680 207.365 109.440 ;
        RECT 207.630 107.825 207.955 108.175 ;
        RECT 210.720 107.825 210.950 107.960 ;
        RECT 211.780 107.825 212.010 107.960 ;
        RECT 207.630 107.645 212.010 107.825 ;
        RECT 207.630 107.070 207.955 107.645 ;
        RECT 210.720 107.500 210.950 107.645 ;
        RECT 211.780 107.500 212.010 107.645 ;
        RECT 211.155 107.340 211.575 107.450 ;
        RECT 211.140 107.150 212.030 107.340 ;
        RECT 207.040 105.450 207.460 105.680 ;
        RECT 203.650 105.380 203.880 105.400 ;
        RECT 203.510 105.270 203.880 105.380 ;
        RECT 204.620 105.270 204.850 105.400 ;
        RECT 203.510 105.090 204.850 105.270 ;
        RECT 203.510 104.940 203.880 105.090 ;
        RECT 204.620 104.940 204.850 105.090 ;
        RECT 206.650 105.260 206.880 105.400 ;
        RECT 207.620 105.260 207.850 105.400 ;
        RECT 206.650 105.070 207.850 105.260 ;
        RECT 206.650 104.940 206.880 105.070 ;
        RECT 207.620 104.940 207.850 105.070 ;
        RECT 203.510 104.740 203.710 104.940 ;
        RECT 204.040 104.740 204.460 104.890 ;
        RECT 207.040 104.740 207.460 104.890 ;
        RECT 203.510 104.520 207.500 104.740 ;
        RECT 203.510 102.620 203.710 104.520 ;
        RECT 207.660 104.350 207.840 104.940 ;
        RECT 211.840 104.880 212.030 107.150 ;
        RECT 213.625 107.000 213.810 109.440 ;
        RECT 214.840 109.210 217.000 110.390 ;
        RECT 224.840 110.040 227.000 111.220 ;
        RECT 214.840 107.550 217.000 108.730 ;
        RECT 224.840 108.380 227.000 109.560 ;
        RECT 214.870 107.000 216.975 107.020 ;
        RECT 213.625 106.815 216.975 107.000 ;
        RECT 214.845 106.770 216.975 106.815 ;
        RECT 214.845 106.760 215.120 106.770 ;
        RECT 224.840 106.720 227.000 107.900 ;
        RECT 210.720 104.730 210.950 104.880 ;
        RECT 211.780 104.730 212.030 104.880 ;
        RECT 210.720 104.570 212.030 104.730 ;
        RECT 210.720 104.420 210.950 104.570 ;
        RECT 211.780 104.420 212.030 104.570 ;
        RECT 207.600 103.245 207.925 104.350 ;
        RECT 211.155 104.200 211.575 104.370 ;
        RECT 211.840 104.200 212.030 104.420 ;
        RECT 208.425 103.970 212.030 104.200 ;
        RECT 206.270 102.800 207.490 103.020 ;
        RECT 203.510 102.470 203.880 102.620 ;
        RECT 204.620 102.470 204.850 102.620 ;
        RECT 203.510 102.290 204.850 102.470 ;
        RECT 203.510 102.160 203.880 102.290 ;
        RECT 204.620 102.160 204.850 102.290 ;
        RECT 203.510 99.840 203.710 102.160 ;
        RECT 204.040 101.940 204.460 102.110 ;
        RECT 206.270 101.940 206.490 102.800 ;
        RECT 207.040 102.670 207.460 102.800 ;
        RECT 207.660 102.620 207.840 103.245 ;
        RECT 206.650 102.500 206.880 102.620 ;
        RECT 207.620 102.500 207.850 102.620 ;
        RECT 206.650 102.310 207.850 102.500 ;
        RECT 206.650 102.160 206.880 102.310 ;
        RECT 207.620 102.160 207.850 102.310 ;
        RECT 204.040 101.720 206.490 101.940 ;
        RECT 207.040 101.960 207.460 102.110 ;
        RECT 208.425 101.960 208.655 103.970 ;
        RECT 207.040 101.880 208.655 101.960 ;
        RECT 207.050 101.730 208.655 101.880 ;
        RECT 211.840 101.800 212.030 103.970 ;
        RECT 210.720 101.675 210.950 101.800 ;
        RECT 211.780 101.675 212.030 101.800 ;
        RECT 214.835 101.680 216.995 102.860 ;
        RECT 224.835 102.510 226.995 103.690 ;
        RECT 210.720 101.515 212.030 101.675 ;
        RECT 210.720 101.340 210.950 101.515 ;
        RECT 211.780 101.340 212.030 101.515 ;
        RECT 211.840 101.335 212.030 101.340 ;
        RECT 211.155 101.060 211.575 101.290 ;
        RECT 206.280 100.030 207.470 100.250 ;
        RECT 203.510 99.690 203.880 99.840 ;
        RECT 204.620 99.690 204.850 99.840 ;
        RECT 203.510 99.510 204.850 99.690 ;
        RECT 203.510 99.380 203.880 99.510 ;
        RECT 204.620 99.380 204.850 99.510 ;
        RECT 203.510 98.295 203.710 99.380 ;
        RECT 204.040 99.170 204.460 99.330 ;
        RECT 206.280 99.170 206.500 100.030 ;
        RECT 207.040 99.890 207.460 100.030 ;
        RECT 207.040 99.205 207.460 99.330 ;
        RECT 204.030 98.950 206.500 99.170 ;
        RECT 207.025 99.100 207.460 99.205 ;
        RECT 207.025 98.995 207.440 99.100 ;
        RECT 211.275 99.000 211.455 101.060 ;
        RECT 214.835 100.020 216.995 101.200 ;
        RECT 224.835 100.850 226.995 102.030 ;
        RECT 203.510 98.095 204.345 98.295 ;
        RECT 204.145 97.340 204.345 98.095 ;
        RECT 207.230 98.075 207.440 98.995 ;
        RECT 211.155 98.770 211.575 99.000 ;
        RECT 214.835 98.360 216.995 99.540 ;
        RECT 224.835 99.190 226.995 100.370 ;
        RECT 211.155 98.075 211.575 98.210 ;
        RECT 207.230 97.865 211.585 98.075 ;
        RECT 207.230 97.860 207.440 97.865 ;
        RECT 204.040 97.110 204.460 97.340 ;
        RECT 203.650 96.900 203.880 97.060 ;
        RECT 204.620 96.940 204.850 97.060 ;
        RECT 204.620 96.900 204.920 96.940 ;
        RECT 203.650 96.730 204.930 96.900 ;
        RECT 203.650 96.600 203.880 96.730 ;
        RECT 204.620 96.600 204.920 96.730 ;
        RECT 204.730 95.960 204.920 96.600 ;
        RECT 204.660 94.855 204.985 95.960 ;
        RECT 208.660 95.480 208.845 97.865 ;
        RECT 214.835 96.700 216.995 97.880 ;
        RECT 224.835 97.530 226.995 98.710 ;
        RECT 210.720 95.480 210.950 95.640 ;
        RECT 211.780 95.480 212.010 95.640 ;
        RECT 208.660 95.295 212.010 95.480 ;
        RECT 204.730 94.280 204.920 94.855 ;
        RECT 203.650 94.135 203.880 94.280 ;
        RECT 204.620 94.135 204.920 94.280 ;
        RECT 206.650 94.150 206.880 94.280 ;
        RECT 203.650 93.965 204.920 94.135 ;
        RECT 203.650 93.820 203.880 93.965 ;
        RECT 204.620 93.820 204.920 93.965 ;
        RECT 205.635 94.125 206.880 94.150 ;
        RECT 207.620 94.125 207.850 94.280 ;
        RECT 208.660 94.125 208.845 95.295 ;
        RECT 210.720 95.180 210.950 95.295 ;
        RECT 211.780 95.180 212.010 95.295 ;
        RECT 211.155 95.015 211.575 95.130 ;
        RECT 214.835 95.040 216.995 96.220 ;
        RECT 224.835 95.870 226.995 97.050 ;
        RECT 205.635 93.940 208.845 94.125 ;
        RECT 209.130 94.830 211.585 95.015 ;
        RECT 205.635 93.935 206.880 93.940 ;
        RECT 204.040 93.605 204.460 93.770 ;
        RECT 205.635 93.605 205.850 93.935 ;
        RECT 206.650 93.820 206.880 93.935 ;
        RECT 207.620 93.820 207.850 93.940 ;
        RECT 207.040 93.610 207.460 93.770 ;
        RECT 209.130 93.610 209.315 94.830 ;
        RECT 204.015 93.390 205.850 93.605 ;
        RECT 207.025 93.425 209.315 93.610 ;
        RECT 209.110 92.385 209.290 93.425 ;
        RECT 214.835 93.380 216.995 94.560 ;
        RECT 224.835 94.210 226.995 95.390 ;
        RECT 210.720 92.385 210.950 92.560 ;
        RECT 211.780 92.385 212.010 92.560 ;
        RECT 209.110 92.205 212.010 92.385 ;
        RECT 203.650 91.380 203.880 91.500 ;
        RECT 204.620 91.450 204.850 91.500 ;
        RECT 204.620 91.380 204.990 91.450 ;
        RECT 203.650 91.190 204.990 91.380 ;
        RECT 206.650 91.360 206.880 91.500 ;
        RECT 207.620 91.360 207.850 91.500 ;
        RECT 209.110 91.360 209.290 92.205 ;
        RECT 210.720 92.100 210.950 92.205 ;
        RECT 211.780 92.100 212.010 92.205 ;
        RECT 211.155 91.885 211.575 92.050 ;
        RECT 212.245 91.885 212.570 92.685 ;
        RECT 203.650 91.040 203.880 91.190 ;
        RECT 204.620 91.040 204.990 91.190 ;
        RECT 204.040 90.825 204.460 90.990 ;
        RECT 203.320 90.760 204.460 90.825 ;
        RECT 203.320 90.410 204.455 90.760 ;
        RECT 203.320 89.300 203.515 90.410 ;
        RECT 203.320 89.000 204.445 89.300 ;
        RECT 203.320 88.885 204.460 89.000 ;
        RECT 203.320 86.590 203.510 88.885 ;
        RECT 204.040 88.770 204.460 88.885 ;
        RECT 204.770 88.720 204.990 91.040 ;
        RECT 206.635 91.180 209.290 91.360 ;
        RECT 209.720 91.685 212.570 91.885 ;
        RECT 214.835 91.720 216.995 92.900 ;
        RECT 224.835 92.550 226.995 93.730 ;
        RECT 206.635 91.040 206.880 91.180 ;
        RECT 207.620 91.040 207.850 91.180 ;
        RECT 206.635 90.060 206.815 91.040 ;
        RECT 207.040 90.835 207.460 90.990 ;
        RECT 209.720 90.835 209.920 91.685 ;
        RECT 212.245 91.580 212.570 91.685 ;
        RECT 207.035 90.635 209.920 90.835 ;
        RECT 214.835 90.060 216.995 91.240 ;
        RECT 224.835 90.890 226.995 92.070 ;
        RECT 206.635 89.880 207.880 90.060 ;
        RECT 207.700 88.720 207.880 89.880 ;
        RECT 210.720 89.335 210.950 89.480 ;
        RECT 211.780 89.335 212.010 89.480 ;
        RECT 203.650 88.575 203.880 88.720 ;
        RECT 204.620 88.575 204.990 88.720 ;
        RECT 203.650 88.385 204.990 88.575 ;
        RECT 203.650 88.260 203.880 88.385 ;
        RECT 204.620 88.260 204.990 88.385 ;
        RECT 206.650 88.570 206.880 88.720 ;
        RECT 207.620 88.570 207.880 88.720 ;
        RECT 209.115 89.175 212.010 89.335 ;
        RECT 209.115 88.570 209.275 89.175 ;
        RECT 210.720 89.020 210.950 89.175 ;
        RECT 211.780 89.020 212.010 89.175 ;
        RECT 211.155 88.790 211.575 88.970 ;
        RECT 206.650 88.410 209.275 88.570 ;
        RECT 209.565 88.610 213.165 88.790 ;
        RECT 206.650 88.260 206.880 88.410 ;
        RECT 207.620 88.405 207.880 88.410 ;
        RECT 207.620 88.260 207.850 88.405 ;
        RECT 204.770 88.240 204.990 88.260 ;
        RECT 204.040 87.980 204.460 88.210 ;
        RECT 204.155 87.005 204.355 87.980 ;
        RECT 204.810 87.540 204.970 88.240 ;
        RECT 207.040 88.065 207.460 88.210 ;
        RECT 209.565 88.065 209.745 88.610 ;
        RECT 207.020 87.885 209.745 88.065 ;
        RECT 212.985 88.535 213.165 88.610 ;
        RECT 204.810 87.380 211.295 87.540 ;
        RECT 212.985 87.430 213.310 88.535 ;
        RECT 214.835 88.400 216.995 89.580 ;
        RECT 224.835 89.230 226.995 90.410 ;
        RECT 211.135 87.290 211.295 87.380 ;
        RECT 213.760 87.290 214.085 88.140 ;
        RECT 211.135 87.130 214.085 87.290 ;
        RECT 210.075 87.005 210.400 87.040 ;
        RECT 213.760 87.035 214.085 87.130 ;
        RECT 204.155 86.805 210.445 87.005 ;
        RECT 203.320 86.250 209.640 86.590 ;
        RECT 209.300 85.675 209.640 86.250 ;
        RECT 210.075 85.935 210.400 86.805 ;
        RECT 211.145 86.615 213.985 86.785 ;
        RECT 214.835 86.740 216.995 87.920 ;
        RECT 224.835 87.570 226.995 88.750 ;
        RECT 211.155 86.450 211.575 86.615 ;
        RECT 210.720 86.280 210.950 86.400 ;
        RECT 211.780 86.280 212.010 86.400 ;
        RECT 210.720 86.100 213.465 86.280 ;
        RECT 210.720 85.940 210.950 86.100 ;
        RECT 211.780 85.940 212.010 86.100 ;
        RECT 211.155 85.675 211.575 85.890 ;
        RECT 209.300 85.335 211.585 85.675 ;
        RECT 203.545 82.365 205.705 83.545 ;
        RECT 211.245 83.495 211.585 85.335 ;
        RECT 210.570 83.245 212.675 83.495 ;
        RECT 213.285 80.970 213.465 86.100 ;
        RECT 212.330 80.790 213.465 80.970 ;
        RECT 212.330 79.160 212.510 80.790 ;
        RECT 213.815 80.480 213.985 86.615 ;
        RECT 214.835 85.080 216.995 86.260 ;
        RECT 224.835 85.910 226.995 87.090 ;
        RECT 214.835 83.770 216.995 84.600 ;
        RECT 224.835 84.250 226.995 85.430 ;
        RECT 214.830 83.420 216.995 83.770 ;
        RECT 224.830 83.420 226.995 83.770 ;
        RECT 222.690 82.615 223.720 82.715 ;
        RECT 224.945 82.615 225.165 83.420 ;
        RECT 222.690 82.395 225.165 82.615 ;
        RECT 222.690 82.325 223.720 82.395 ;
        RECT 212.860 80.230 214.965 80.480 ;
        RECT 212.330 78.980 220.090 79.160 ;
        RECT 210.205 78.780 210.530 78.830 ;
        RECT 206.870 77.780 207.870 78.780 ;
        RECT 209.560 77.780 210.560 78.780 ;
        RECT 211.340 78.750 211.665 78.830 ;
        RECT 218.815 78.750 219.140 78.840 ;
        RECT 219.910 78.780 220.090 78.980 ;
        RECT 207.180 76.360 207.420 77.780 ;
        RECT 210.190 77.725 210.530 77.780 ;
        RECT 211.300 77.750 212.300 78.750 ;
        RECT 218.160 77.750 219.160 78.750 ;
        RECT 219.900 77.780 220.900 78.780 ;
        RECT 222.590 77.780 223.590 78.780 ;
        RECT 210.190 77.050 210.520 77.725 ;
        RECT 211.340 77.050 211.670 77.750 ;
        RECT 218.790 77.735 219.140 77.750 ;
        RECT 218.790 77.050 219.120 77.735 ;
        RECT 219.940 77.050 220.270 77.780 ;
        RECT 208.920 76.560 212.680 76.850 ;
        RECT 217.780 76.560 221.540 76.850 ;
        RECT 208.915 76.520 212.685 76.560 ;
        RECT 205.030 76.140 205.260 76.270 ;
        RECT 206.000 76.140 206.230 76.270 ;
        RECT 207.140 76.140 207.470 76.360 ;
        RECT 205.030 75.940 207.470 76.140 ;
        RECT 205.030 75.810 205.260 75.940 ;
        RECT 206.000 75.810 206.230 75.940 ;
        RECT 207.140 75.770 207.470 75.940 ;
        RECT 208.430 76.120 208.760 76.350 ;
        RECT 208.915 76.330 209.335 76.520 ;
        RECT 212.265 76.330 212.685 76.520 ;
        RECT 217.775 76.520 221.545 76.560 ;
        RECT 217.775 76.330 218.195 76.520 ;
        RECT 221.125 76.330 221.545 76.520 ;
        RECT 223.040 76.360 223.280 77.780 ;
        RECT 209.540 76.120 209.770 76.280 ;
        RECT 211.830 76.190 212.060 76.280 ;
        RECT 212.890 76.190 213.120 76.280 ;
        RECT 208.430 75.910 209.850 76.120 ;
        RECT 211.330 75.930 213.120 76.190 ;
        RECT 208.430 75.760 208.760 75.910 ;
        RECT 209.540 75.820 209.770 75.910 ;
        RECT 205.420 75.570 205.840 75.760 ;
        RECT 208.915 75.570 209.335 75.770 ;
        RECT 211.330 75.640 211.590 75.930 ;
        RECT 211.830 75.820 212.060 75.930 ;
        RECT 212.890 75.820 213.120 75.930 ;
        RECT 217.340 76.190 217.570 76.280 ;
        RECT 218.400 76.190 218.630 76.280 ;
        RECT 217.340 75.930 219.130 76.190 ;
        RECT 220.690 76.120 220.920 76.280 ;
        RECT 221.700 76.120 222.030 76.350 ;
        RECT 217.340 75.820 217.570 75.930 ;
        RECT 218.400 75.820 218.630 75.930 ;
        RECT 218.870 75.640 219.130 75.930 ;
        RECT 220.610 75.910 222.030 76.120 ;
        RECT 220.690 75.820 220.920 75.910 ;
        RECT 209.520 75.570 209.850 75.640 ;
        RECT 211.300 75.570 211.630 75.640 ;
        RECT 205.380 75.310 211.630 75.570 ;
        RECT 209.520 75.050 209.850 75.310 ;
        RECT 211.300 75.050 211.630 75.310 ;
        RECT 218.830 75.570 219.160 75.640 ;
        RECT 220.610 75.570 220.940 75.640 ;
        RECT 221.125 75.570 221.545 75.770 ;
        RECT 221.700 75.760 222.030 75.910 ;
        RECT 222.990 76.140 223.320 76.360 ;
        RECT 224.230 76.140 224.460 76.270 ;
        RECT 225.200 76.140 225.430 76.270 ;
        RECT 222.990 75.940 225.430 76.140 ;
        RECT 222.990 75.770 223.320 75.940 ;
        RECT 224.230 75.810 224.460 75.940 ;
        RECT 225.200 75.810 225.430 75.940 ;
        RECT 224.620 75.570 225.040 75.760 ;
        RECT 218.830 75.310 225.080 75.570 ;
        RECT 218.830 75.050 219.160 75.310 ;
        RECT 220.610 75.050 220.940 75.310 ;
        RECT 208.430 73.720 208.760 74.000 ;
        RECT 210.180 73.720 210.510 73.990 ;
        RECT 219.950 73.720 220.280 73.990 ;
        RECT 221.700 73.720 222.030 74.000 ;
        RECT 205.400 73.460 211.600 73.720 ;
        RECT 205.410 73.290 205.830 73.460 ;
        RECT 208.430 73.410 208.760 73.460 ;
        RECT 208.925 73.280 209.345 73.460 ;
        RECT 210.180 73.400 210.510 73.460 ;
        RECT 208.490 73.120 208.720 73.230 ;
        RECT 209.530 73.120 209.860 73.300 ;
        RECT 208.490 72.910 209.860 73.120 ;
        RECT 208.490 72.770 208.720 72.910 ;
        RECT 208.925 72.510 209.345 72.720 ;
        RECT 209.530 72.710 209.860 72.910 ;
        RECT 211.340 73.100 211.600 73.460 ;
        RECT 218.860 73.460 225.060 73.720 ;
        RECT 211.830 73.100 212.060 73.200 ;
        RECT 212.890 73.100 213.120 73.200 ;
        RECT 211.340 72.840 213.120 73.100 ;
        RECT 211.830 72.740 212.060 72.840 ;
        RECT 212.890 72.740 213.120 72.840 ;
        RECT 217.340 73.100 217.570 73.200 ;
        RECT 218.400 73.100 218.630 73.200 ;
        RECT 218.860 73.100 219.120 73.460 ;
        RECT 219.950 73.400 220.280 73.460 ;
        RECT 217.340 72.840 219.120 73.100 ;
        RECT 220.600 73.120 220.930 73.300 ;
        RECT 221.115 73.280 221.535 73.460 ;
        RECT 221.700 73.410 222.030 73.460 ;
        RECT 224.630 73.290 225.050 73.460 ;
        RECT 221.740 73.120 221.970 73.230 ;
        RECT 220.600 72.910 221.970 73.120 ;
        RECT 217.340 72.740 217.570 72.840 ;
        RECT 218.400 72.740 218.630 72.840 ;
        RECT 220.600 72.710 220.930 72.910 ;
        RECT 221.740 72.770 221.970 72.910 ;
        RECT 212.265 72.510 212.685 72.690 ;
        RECT 208.920 72.460 212.685 72.510 ;
        RECT 217.775 72.510 218.195 72.690 ;
        RECT 221.115 72.510 221.535 72.720 ;
        RECT 217.775 72.460 221.540 72.510 ;
        RECT 208.920 72.180 212.680 72.460 ;
        RECT 217.780 72.180 221.540 72.460 ;
        RECT 207.140 65.230 207.470 65.720 ;
        RECT 213.900 65.510 214.190 65.550 ;
        RECT 215.010 65.510 215.335 66.365 ;
        RECT 213.900 65.320 215.755 65.510 ;
        RECT 213.995 65.315 215.755 65.320 ;
        RECT 215.010 65.260 215.335 65.315 ;
        RECT 207.110 65.070 210.960 65.230 ;
        RECT 206.740 65.020 210.960 65.070 ;
        RECT 215.560 65.130 215.755 65.315 ;
        RECT 222.990 65.230 223.320 65.720 ;
        RECT 206.740 64.840 207.740 65.020 ;
        RECT 209.930 64.840 210.930 65.020 ;
        RECT 215.560 64.935 216.575 65.130 ;
        RECT 219.500 65.070 223.350 65.230 ;
        RECT 219.500 65.020 223.720 65.070 ;
        RECT 216.270 64.875 216.560 64.935 ;
        RECT 219.530 64.840 220.530 65.020 ;
        RECT 222.720 64.840 223.720 65.020 ;
      LAYER via ;
        RECT 213.925 113.520 214.185 113.780 ;
        RECT 213.925 113.200 214.185 113.460 ;
        RECT 213.925 112.880 214.185 113.140 ;
        RECT 207.660 107.815 207.920 108.075 ;
        RECT 207.660 107.495 207.920 107.755 ;
        RECT 207.660 107.175 207.920 107.435 ;
        RECT 207.630 103.990 207.890 104.250 ;
        RECT 207.630 103.670 207.890 103.930 ;
        RECT 207.630 103.350 207.890 103.610 ;
        RECT 204.690 95.600 204.950 95.860 ;
        RECT 204.690 95.280 204.950 95.540 ;
        RECT 204.690 94.960 204.950 95.220 ;
        RECT 212.275 92.325 212.535 92.585 ;
        RECT 212.275 92.005 212.535 92.265 ;
        RECT 212.275 91.685 212.535 91.945 ;
        RECT 213.015 88.175 213.275 88.435 ;
        RECT 213.015 87.855 213.275 88.115 ;
        RECT 213.015 87.535 213.275 87.795 ;
        RECT 213.790 87.780 214.050 88.040 ;
        RECT 213.790 87.460 214.050 87.720 ;
        RECT 213.790 87.140 214.050 87.400 ;
        RECT 210.105 86.680 210.365 86.940 ;
        RECT 210.105 86.360 210.365 86.620 ;
        RECT 210.105 86.040 210.365 86.300 ;
        RECT 222.755 82.390 223.015 82.650 ;
        RECT 223.075 82.390 223.335 82.650 ;
        RECT 223.395 82.390 223.655 82.650 ;
        RECT 210.235 78.470 210.495 78.730 ;
        RECT 210.235 78.150 210.495 78.410 ;
        RECT 210.235 77.830 210.495 78.090 ;
        RECT 211.370 78.470 211.630 78.730 ;
        RECT 211.370 78.150 211.630 78.410 ;
        RECT 211.370 77.830 211.630 78.090 ;
        RECT 218.845 78.480 219.105 78.740 ;
        RECT 218.845 78.160 219.105 78.420 ;
        RECT 218.845 77.840 219.105 78.100 ;
        RECT 210.225 77.215 210.485 77.475 ;
        RECT 211.375 77.215 211.635 77.475 ;
        RECT 218.825 77.215 219.085 77.475 ;
        RECT 219.975 77.215 220.235 77.475 ;
        RECT 207.175 75.935 207.435 76.195 ;
        RECT 208.465 75.925 208.725 76.185 ;
        RECT 221.735 75.925 221.995 76.185 ;
        RECT 209.555 75.215 209.815 75.475 ;
        RECT 211.335 75.215 211.595 75.475 ;
        RECT 223.025 75.935 223.285 76.195 ;
        RECT 218.865 75.215 219.125 75.475 ;
        RECT 220.645 75.215 220.905 75.475 ;
        RECT 208.465 73.575 208.725 73.835 ;
        RECT 210.215 73.565 210.475 73.825 ;
        RECT 209.565 72.875 209.825 73.135 ;
        RECT 219.985 73.565 220.245 73.825 ;
        RECT 221.735 73.575 221.995 73.835 ;
        RECT 220.635 72.875 220.895 73.135 ;
        RECT 215.040 66.005 215.300 66.265 ;
        RECT 207.175 65.295 207.435 65.555 ;
        RECT 215.040 65.685 215.300 65.945 ;
        RECT 215.040 65.365 215.300 65.625 ;
        RECT 223.025 65.295 223.285 65.555 ;
      LAYER met2 ;
        RECT 213.845 112.825 214.270 113.830 ;
        RECT 207.580 107.120 208.005 108.125 ;
        RECT 207.655 104.300 207.905 107.120 ;
        RECT 207.550 103.295 207.975 104.300 ;
        RECT 204.610 94.905 205.035 95.910 ;
        RECT 204.700 80.265 204.950 94.905 ;
        RECT 207.655 80.885 207.905 103.295 ;
        RECT 213.955 97.980 214.155 112.825 ;
        RECT 212.305 97.780 214.155 97.980 ;
        RECT 212.305 92.635 212.505 97.780 ;
        RECT 212.195 91.630 212.620 92.635 ;
        RECT 212.305 88.890 212.505 91.630 ;
        RECT 212.305 88.690 214.675 88.890 ;
        RECT 210.025 86.960 210.450 86.990 ;
        RECT 212.305 86.960 212.505 88.690 ;
        RECT 212.935 87.480 213.360 88.485 ;
        RECT 213.710 87.865 214.140 88.090 ;
        RECT 210.025 86.760 212.505 86.960 ;
        RECT 210.025 85.985 210.450 86.760 ;
        RECT 213.040 86.000 213.260 87.480 ;
        RECT 213.710 87.085 214.135 87.865 ;
        RECT 213.040 85.780 213.460 86.000 ;
        RECT 207.655 80.635 211.635 80.885 ;
        RECT 204.700 80.015 210.520 80.265 ;
        RECT 210.270 78.780 210.520 80.015 ;
        RECT 211.385 78.780 211.635 80.635 ;
        RECT 213.240 79.575 213.460 85.780 ;
        RECT 213.870 80.090 214.120 87.085 ;
        RECT 214.475 82.630 214.675 88.690 ;
        RECT 222.640 82.630 223.770 82.665 ;
        RECT 214.475 82.430 223.770 82.630 ;
        RECT 222.640 82.375 223.770 82.430 ;
        RECT 213.870 79.840 219.075 80.090 ;
        RECT 213.240 79.355 215.285 79.575 ;
        RECT 210.155 77.775 210.580 78.780 ;
        RECT 211.290 77.775 211.715 78.780 ;
        RECT 210.270 77.590 210.520 77.775 ;
        RECT 211.385 77.590 211.635 77.775 ;
        RECT 210.140 77.100 210.570 77.590 ;
        RECT 211.290 77.100 211.720 77.590 ;
        RECT 207.090 75.820 207.520 76.310 ;
        RECT 207.170 65.670 207.440 75.820 ;
        RECT 208.380 75.810 208.810 76.300 ;
        RECT 208.480 73.950 208.750 75.810 ;
        RECT 209.550 75.590 209.820 75.660 ;
        RECT 209.470 75.100 209.900 75.590 ;
        RECT 208.380 73.460 208.810 73.950 ;
        RECT 208.480 73.360 208.750 73.460 ;
        RECT 209.550 73.250 209.820 75.100 ;
        RECT 210.200 73.940 210.480 77.100 ;
        RECT 211.360 75.590 211.630 77.100 ;
        RECT 211.250 75.100 211.680 75.590 ;
        RECT 210.130 73.450 210.560 73.940 ;
        RECT 209.480 72.760 209.910 73.250 ;
        RECT 215.065 66.315 215.285 79.355 ;
        RECT 218.825 78.790 219.075 79.840 ;
        RECT 218.765 77.785 219.190 78.790 ;
        RECT 218.825 77.590 219.075 77.785 ;
        RECT 218.740 77.100 219.170 77.590 ;
        RECT 219.890 77.100 220.320 77.590 ;
        RECT 218.830 75.590 219.100 77.100 ;
        RECT 218.780 75.100 219.210 75.590 ;
        RECT 219.980 73.940 220.260 77.100 ;
        RECT 221.650 75.810 222.080 76.300 ;
        RECT 222.940 75.820 223.370 76.310 ;
        RECT 220.640 75.590 220.910 75.660 ;
        RECT 220.560 75.100 220.990 75.590 ;
        RECT 219.900 73.450 220.330 73.940 ;
        RECT 220.640 73.250 220.910 75.100 ;
        RECT 221.710 73.950 221.980 75.810 ;
        RECT 221.650 73.460 222.080 73.950 ;
        RECT 221.710 73.360 221.980 73.460 ;
        RECT 220.550 72.760 220.980 73.250 ;
        RECT 207.090 65.180 207.520 65.670 ;
        RECT 214.960 65.310 215.385 66.315 ;
        RECT 223.020 65.670 223.290 75.820 ;
        RECT 222.940 65.180 223.370 65.670 ;
  END
END sky130_ef_ip__xtal_osc_16M_DI
END LIBRARY

