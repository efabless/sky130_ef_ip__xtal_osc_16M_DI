VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__xtal_osc_16M_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__xtal_osc_16M_DI ;
  ORIGIN 0.000 0.000 ;
  SIZE 454.445 BY 211.800 ;
  PIN dout
    ANTENNADIFFAREA 0.435000 ;
    PORT
      LAYER met2 ;
        RECT 142.785 -3.280 143.065 60.465 ;
    END
  END dout
  PIN in
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.526800 ;
    PORT
      LAYER met2 ;
        RECT 448.925 134.970 449.565 218.525 ;
    END
  END in
  PIN ena
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER met2 ;
        RECT 137.535 -3.280 137.815 61.955 ;
    END
  END ena
  PIN stdby
    ANTENNAGATEAREA 0.510000 ;
    PORT
      LAYER met2 ;
        RECT 150.220 -3.280 150.500 62.785 ;
    END
  END stdby
  PIN out
    PORT
      LAYER met2 ;
        RECT 3.925 134.970 4.565 218.525 ;
    END
  END out
  PIN vssd1
    ANTENNADIFFAREA 21.305099 ;
    PORT
      LAYER met4 ;
        RECT 116.420 0.000 118.020 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.750 0.000 123.350 211.800 ;
    END
  END vssd1
  PIN vdda1
    ANTENNADIFFAREA 98.890800 ;
    PORT
      LAYER met4 ;
        RECT 155.695 0.000 157.295 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.550 0.000 153.150 211.800 ;
    END
  END vdda1
  PIN vccd1
    ANTENNADIFFAREA 4.959600 ;
    PORT
      LAYER met4 ;
        RECT 145.755 0.000 147.355 211.800 ;
    END
  END vccd1
  PIN vssa1
    ANTENNADIFFAREA 81.684601 ;
    PORT
      LAYER met4 ;
        RECT 135.235 0.000 136.835 211.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 130.710 0.000 132.310 211.800 ;
    END
  END vssa1
  OBS
      LAYER li1 ;
        RECT 130.565 62.550 158.160 116.595 ;
      LAYER met1 ;
        RECT 114.890 60.240 158.190 117.060 ;
      LAYER met2 ;
        RECT 4.845 134.690 448.645 135.970 ;
        RECT 4.565 63.065 448.925 134.690 ;
        RECT 4.565 62.235 149.940 63.065 ;
        RECT 4.565 0.000 137.255 62.235 ;
        RECT 138.095 60.745 149.940 62.235 ;
        RECT 138.095 0.000 142.505 60.745 ;
        RECT 143.345 0.000 149.940 60.745 ;
        RECT 150.780 0.000 448.925 63.065 ;
      LAYER met3 ;
        RECT 116.020 62.420 158.420 117.060 ;
  END
END sky130_ef_ip__xtal_osc_16M_DI
END LIBRARY

