magic
tech sky130A
magscale 1 2
timestamp 1528466069
<< checkpaint >>
rect -475 -1916 91173 44965
<< metal1 >>
rect 22978 12693 27085 12704
rect 22978 12513 23294 12693
rect 23602 12690 27085 12693
rect 23602 12513 24359 12690
rect 22978 12510 24359 12513
rect 24667 12510 27085 12690
rect 22978 12508 27085 12510
rect 28557 12209 28757 12708
rect 28557 12093 28608 12209
rect 28724 12093 28757 12209
rect 28557 12048 28757 12093
<< via1 >>
rect 27792 23258 27908 23374
rect 29521 23257 29637 23373
rect 23294 12513 23602 12693
rect 24359 12510 24667 12690
rect 27553 12563 27669 12679
rect 30083 12557 30199 12673
rect 28608 12093 28724 12209
<< metal2 >>
rect 785 27194 913 43705
rect 89785 27194 89913 43705
rect 785 26994 27947 27194
rect 27747 23374 27947 26994
rect 27747 23258 27792 23374
rect 27908 23258 27947 23374
rect 27747 23212 27947 23258
rect 29485 26994 89913 27194
rect 29485 23373 29685 26994
rect 29485 23257 29521 23373
rect 29637 23257 29685 23373
rect 29485 23212 29685 23257
rect 22978 12693 25057 12704
rect 22978 12513 23294 12693
rect 23602 12690 25057 12693
rect 23602 12513 24359 12690
rect 22978 12510 24359 12513
rect 24667 12510 25057 12690
rect 22978 12508 25057 12510
rect 27507 12679 27707 12708
rect 27507 12563 27553 12679
rect 27669 12563 27707 12679
rect 30043 12673 30243 12708
rect 27507 0 27707 12563
rect 30043 12557 30083 12673
rect 30199 12557 30243 12673
rect 28557 12209 28757 12330
rect 28557 12093 28608 12209
rect 28724 12093 28757 12209
rect 28557 0 28757 12093
rect 30043 0 30243 12557
rect 27507 -656 27563 0
rect 28557 -656 28613 0
rect 30044 -656 30100 0
<< via2 >>
rect 26148 23324 26204 23380
rect 26228 23324 26284 23380
rect 26308 23324 26364 23380
rect 26388 23324 26444 23380
rect 27053 23324 27109 23380
rect 27133 23324 27189 23380
rect 27213 23324 27269 23380
rect 27293 23324 27349 23380
rect 26148 23235 26204 23291
rect 26228 23235 26284 23291
rect 26308 23235 26364 23291
rect 26388 23235 26444 23291
rect 27053 23230 27109 23286
rect 27133 23230 27189 23286
rect 27213 23230 27269 23286
rect 27293 23230 27349 23286
rect 30316 23324 30372 23380
rect 30396 23324 30452 23380
rect 30476 23324 30532 23380
rect 30556 23324 30612 23380
rect 31145 23324 31201 23380
rect 31225 23324 31281 23380
rect 31305 23324 31361 23380
rect 31385 23324 31441 23380
rect 23298 12620 23354 12676
rect 23378 12620 23434 12676
rect 23458 12620 23514 12676
rect 23538 12620 23594 12676
rect 23298 12531 23354 12587
rect 23378 12531 23434 12587
rect 23458 12531 23514 12587
rect 23538 12531 23594 12587
rect 24363 12620 24419 12676
rect 24443 12620 24499 12676
rect 24523 12620 24579 12676
rect 24603 12620 24659 12676
rect 24363 12526 24419 12582
rect 24443 12526 24499 12582
rect 24523 12526 24579 12582
rect 24603 12526 24659 12582
rect 29169 12598 29225 12654
rect 29249 12598 29305 12654
rect 29329 12598 29385 12654
rect 29409 12598 29465 12654
rect 29169 12509 29225 12565
rect 29249 12509 29305 12565
rect 29329 12509 29385 12565
rect 29409 12509 29465 12565
<< metal3 >>
rect 26054 23384 27679 23412
rect 26054 23320 26144 23384
rect 26208 23320 26224 23384
rect 26288 23320 26304 23384
rect 26368 23320 26384 23384
rect 26448 23320 27049 23384
rect 27113 23320 27129 23384
rect 27193 23320 27209 23384
rect 27273 23320 27289 23384
rect 27353 23320 27679 23384
rect 26054 23295 27679 23320
rect 26054 23231 26144 23295
rect 26208 23231 26224 23295
rect 26288 23231 26304 23295
rect 26368 23231 26384 23295
rect 26448 23290 27679 23295
rect 26448 23231 27049 23290
rect 26054 23226 27049 23231
rect 27113 23226 27129 23290
rect 27193 23226 27209 23290
rect 27273 23226 27289 23290
rect 27353 23226 27679 23290
rect 30056 23384 31684 23412
rect 30056 23320 30312 23384
rect 30376 23320 30392 23384
rect 30456 23320 30472 23384
rect 30536 23320 30552 23384
rect 30616 23320 31141 23384
rect 31205 23320 31221 23384
rect 31285 23320 31301 23384
rect 31365 23320 31381 23384
rect 31445 23320 31684 23384
rect 30056 23287 31684 23320
rect 26054 23210 27679 23226
rect 23204 12680 24829 12708
rect 23204 12616 23294 12680
rect 23358 12616 23374 12680
rect 23438 12616 23454 12680
rect 23518 12616 23534 12680
rect 23598 12616 24359 12680
rect 24423 12616 24439 12680
rect 24503 12616 24519 12680
rect 24583 12616 24599 12680
rect 24663 12616 24829 12680
rect 23204 12591 24829 12616
rect 23204 12527 23294 12591
rect 23358 12527 23374 12591
rect 23438 12527 23454 12591
rect 23518 12527 23534 12591
rect 23598 12586 24829 12591
rect 23598 12527 24359 12586
rect 23204 12522 24359 12527
rect 24423 12522 24439 12586
rect 24503 12522 24519 12586
rect 24583 12522 24599 12586
rect 24663 12522 24829 12586
rect 23204 12506 24829 12522
rect 29075 12658 29659 12686
rect 29075 12594 29165 12658
rect 29229 12594 29245 12658
rect 29309 12594 29325 12658
rect 29389 12594 29405 12658
rect 29469 12594 29659 12658
rect 29075 12569 29659 12594
rect 29075 12505 29165 12569
rect 29229 12505 29245 12569
rect 29309 12505 29325 12569
rect 29389 12505 29405 12569
rect 29469 12505 29659 12569
rect 29075 12484 29659 12505
<< via3 >>
rect 26144 23380 26208 23384
rect 26144 23324 26148 23380
rect 26148 23324 26204 23380
rect 26204 23324 26208 23380
rect 26144 23320 26208 23324
rect 26224 23380 26288 23384
rect 26224 23324 26228 23380
rect 26228 23324 26284 23380
rect 26284 23324 26288 23380
rect 26224 23320 26288 23324
rect 26304 23380 26368 23384
rect 26304 23324 26308 23380
rect 26308 23324 26364 23380
rect 26364 23324 26368 23380
rect 26304 23320 26368 23324
rect 26384 23380 26448 23384
rect 26384 23324 26388 23380
rect 26388 23324 26444 23380
rect 26444 23324 26448 23380
rect 26384 23320 26448 23324
rect 27049 23380 27113 23384
rect 27049 23324 27053 23380
rect 27053 23324 27109 23380
rect 27109 23324 27113 23380
rect 27049 23320 27113 23324
rect 27129 23380 27193 23384
rect 27129 23324 27133 23380
rect 27133 23324 27189 23380
rect 27189 23324 27193 23380
rect 27129 23320 27193 23324
rect 27209 23380 27273 23384
rect 27209 23324 27213 23380
rect 27213 23324 27269 23380
rect 27269 23324 27273 23380
rect 27209 23320 27273 23324
rect 27289 23380 27353 23384
rect 27289 23324 27293 23380
rect 27293 23324 27349 23380
rect 27349 23324 27353 23380
rect 27289 23320 27353 23324
rect 26144 23291 26208 23295
rect 26144 23235 26148 23291
rect 26148 23235 26204 23291
rect 26204 23235 26208 23291
rect 26144 23231 26208 23235
rect 26224 23291 26288 23295
rect 26224 23235 26228 23291
rect 26228 23235 26284 23291
rect 26284 23235 26288 23291
rect 26224 23231 26288 23235
rect 26304 23291 26368 23295
rect 26304 23235 26308 23291
rect 26308 23235 26364 23291
rect 26364 23235 26368 23291
rect 26304 23231 26368 23235
rect 26384 23291 26448 23295
rect 26384 23235 26388 23291
rect 26388 23235 26444 23291
rect 26444 23235 26448 23291
rect 26384 23231 26448 23235
rect 27049 23286 27113 23290
rect 27049 23230 27053 23286
rect 27053 23230 27109 23286
rect 27109 23230 27113 23286
rect 27049 23226 27113 23230
rect 27129 23286 27193 23290
rect 27129 23230 27133 23286
rect 27133 23230 27189 23286
rect 27189 23230 27193 23286
rect 27129 23226 27193 23230
rect 27209 23286 27273 23290
rect 27209 23230 27213 23286
rect 27213 23230 27269 23286
rect 27269 23230 27273 23286
rect 27209 23226 27273 23230
rect 27289 23286 27353 23290
rect 27289 23230 27293 23286
rect 27293 23230 27349 23286
rect 27349 23230 27353 23286
rect 27289 23226 27353 23230
rect 30312 23380 30376 23384
rect 30312 23324 30316 23380
rect 30316 23324 30372 23380
rect 30372 23324 30376 23380
rect 30312 23320 30376 23324
rect 30392 23380 30456 23384
rect 30392 23324 30396 23380
rect 30396 23324 30452 23380
rect 30452 23324 30456 23380
rect 30392 23320 30456 23324
rect 30472 23380 30536 23384
rect 30472 23324 30476 23380
rect 30476 23324 30532 23380
rect 30532 23324 30536 23380
rect 30472 23320 30536 23324
rect 30552 23380 30616 23384
rect 30552 23324 30556 23380
rect 30556 23324 30612 23380
rect 30612 23324 30616 23380
rect 30552 23320 30616 23324
rect 31141 23380 31205 23384
rect 31141 23324 31145 23380
rect 31145 23324 31201 23380
rect 31201 23324 31205 23380
rect 31141 23320 31205 23324
rect 31221 23380 31285 23384
rect 31221 23324 31225 23380
rect 31225 23324 31281 23380
rect 31281 23324 31285 23380
rect 31221 23320 31285 23324
rect 31301 23380 31365 23384
rect 31301 23324 31305 23380
rect 31305 23324 31361 23380
rect 31361 23324 31365 23380
rect 31301 23320 31365 23324
rect 31381 23380 31445 23384
rect 31381 23324 31385 23380
rect 31385 23324 31441 23380
rect 31441 23324 31445 23380
rect 31381 23320 31445 23324
rect 23294 12676 23358 12680
rect 23294 12620 23298 12676
rect 23298 12620 23354 12676
rect 23354 12620 23358 12676
rect 23294 12616 23358 12620
rect 23374 12676 23438 12680
rect 23374 12620 23378 12676
rect 23378 12620 23434 12676
rect 23434 12620 23438 12676
rect 23374 12616 23438 12620
rect 23454 12676 23518 12680
rect 23454 12620 23458 12676
rect 23458 12620 23514 12676
rect 23514 12620 23518 12676
rect 23454 12616 23518 12620
rect 23534 12676 23598 12680
rect 23534 12620 23538 12676
rect 23538 12620 23594 12676
rect 23594 12620 23598 12676
rect 23534 12616 23598 12620
rect 24359 12676 24423 12680
rect 24359 12620 24363 12676
rect 24363 12620 24419 12676
rect 24419 12620 24423 12676
rect 24359 12616 24423 12620
rect 24439 12676 24503 12680
rect 24439 12620 24443 12676
rect 24443 12620 24499 12676
rect 24499 12620 24503 12676
rect 24439 12616 24503 12620
rect 24519 12676 24583 12680
rect 24519 12620 24523 12676
rect 24523 12620 24579 12676
rect 24579 12620 24583 12676
rect 24519 12616 24583 12620
rect 24599 12676 24663 12680
rect 24599 12620 24603 12676
rect 24603 12620 24659 12676
rect 24659 12620 24663 12676
rect 24599 12616 24663 12620
rect 23294 12587 23358 12591
rect 23294 12531 23298 12587
rect 23298 12531 23354 12587
rect 23354 12531 23358 12587
rect 23294 12527 23358 12531
rect 23374 12587 23438 12591
rect 23374 12531 23378 12587
rect 23378 12531 23434 12587
rect 23434 12531 23438 12587
rect 23374 12527 23438 12531
rect 23454 12587 23518 12591
rect 23454 12531 23458 12587
rect 23458 12531 23514 12587
rect 23514 12531 23518 12587
rect 23454 12527 23518 12531
rect 23534 12587 23598 12591
rect 23534 12531 23538 12587
rect 23538 12531 23594 12587
rect 23594 12531 23598 12587
rect 23534 12527 23598 12531
rect 24359 12582 24423 12586
rect 24359 12526 24363 12582
rect 24363 12526 24419 12582
rect 24419 12526 24423 12582
rect 24359 12522 24423 12526
rect 24439 12582 24503 12586
rect 24439 12526 24443 12582
rect 24443 12526 24499 12582
rect 24499 12526 24503 12582
rect 24439 12522 24503 12526
rect 24519 12582 24583 12586
rect 24519 12526 24523 12582
rect 24523 12526 24579 12582
rect 24579 12526 24583 12582
rect 24519 12522 24583 12526
rect 24599 12582 24663 12586
rect 24599 12526 24603 12582
rect 24603 12526 24659 12582
rect 24659 12526 24663 12582
rect 24599 12522 24663 12526
rect 29165 12654 29229 12658
rect 29165 12598 29169 12654
rect 29169 12598 29225 12654
rect 29225 12598 29229 12654
rect 29165 12594 29229 12598
rect 29245 12654 29309 12658
rect 29245 12598 29249 12654
rect 29249 12598 29305 12654
rect 29305 12598 29309 12654
rect 29245 12594 29309 12598
rect 29325 12654 29389 12658
rect 29325 12598 29329 12654
rect 29329 12598 29385 12654
rect 29385 12598 29389 12654
rect 29325 12594 29389 12598
rect 29405 12654 29469 12658
rect 29405 12598 29409 12654
rect 29409 12598 29465 12654
rect 29465 12598 29469 12654
rect 29405 12594 29469 12598
rect 29165 12565 29229 12569
rect 29165 12509 29169 12565
rect 29169 12509 29225 12565
rect 29225 12509 29229 12565
rect 29165 12505 29229 12509
rect 29245 12565 29309 12569
rect 29245 12509 29249 12565
rect 29249 12509 29305 12565
rect 29305 12509 29309 12565
rect 29245 12505 29309 12509
rect 29325 12565 29389 12569
rect 29325 12509 29329 12565
rect 29329 12509 29385 12565
rect 29385 12509 29389 12565
rect 29325 12505 29389 12509
rect 29405 12565 29469 12569
rect 29405 12509 29409 12565
rect 29409 12509 29465 12565
rect 29465 12509 29469 12565
rect 29405 12505 29469 12509
<< metal4 >>
rect 23284 12680 23604 42360
rect 23284 12616 23294 12680
rect 23358 12616 23374 12680
rect 23438 12616 23454 12680
rect 23518 12616 23534 12680
rect 23598 12616 23604 12680
rect 23284 12591 23604 12616
rect 23284 12527 23294 12591
rect 23358 12527 23374 12591
rect 23438 12527 23454 12591
rect 23518 12527 23534 12591
rect 23598 12527 23604 12591
rect 23284 0 23604 12527
rect 24350 12680 24670 42360
rect 24350 12616 24359 12680
rect 24423 12616 24439 12680
rect 24503 12616 24519 12680
rect 24583 12616 24599 12680
rect 24663 12616 24670 12680
rect 24350 12586 24670 12616
rect 24350 12522 24359 12586
rect 24423 12522 24439 12586
rect 24503 12522 24519 12586
rect 24583 12522 24599 12586
rect 24663 12522 24670 12586
rect 24350 0 24670 12522
rect 26142 23384 26462 42360
rect 26142 23320 26144 23384
rect 26208 23320 26224 23384
rect 26288 23320 26304 23384
rect 26368 23320 26384 23384
rect 26448 23320 26462 23384
rect 26142 23295 26462 23320
rect 26142 23231 26144 23295
rect 26208 23231 26224 23295
rect 26288 23231 26304 23295
rect 26368 23231 26384 23295
rect 26448 23231 26462 23295
rect 26142 0 26462 23231
rect 27047 23384 27367 42360
rect 27047 23320 27049 23384
rect 27113 23320 27129 23384
rect 27193 23320 27209 23384
rect 27273 23320 27289 23384
rect 27353 23320 27367 23384
rect 27047 23290 27367 23320
rect 27047 23226 27049 23290
rect 27113 23226 27129 23290
rect 27193 23226 27209 23290
rect 27273 23226 27289 23290
rect 27353 23226 27367 23290
rect 27047 0 27367 23226
rect 29151 12658 29471 42360
rect 29151 12594 29165 12658
rect 29229 12594 29245 12658
rect 29309 12594 29325 12658
rect 29389 12594 29405 12658
rect 29469 12594 29471 12658
rect 29151 12569 29471 12594
rect 29151 12505 29165 12569
rect 29229 12505 29245 12569
rect 29309 12505 29325 12569
rect 29389 12505 29405 12569
rect 29469 12505 29471 12569
rect 29151 0 29471 12505
rect 30310 23384 30630 42360
rect 30310 23320 30312 23384
rect 30376 23320 30392 23384
rect 30456 23320 30472 23384
rect 30536 23320 30552 23384
rect 30616 23320 30630 23384
rect 30310 0 30630 23320
rect 31139 23384 31459 42360
rect 31139 23320 31141 23384
rect 31205 23320 31221 23384
rect 31285 23320 31301 23384
rect 31365 23320 31381 23384
rect 31445 23320 31459 23384
rect 31139 0 31459 23320
use sky130_ef_ip__xtal_osc_16M  sky130_ef_ip__xtal_osc_16M_0
timestamp 1528466069
transform 0 1 28469 -1 0 25872
box 2460 -2440 13388 3256
<< labels >>
flabel metal2 s 785 42249 913 43705 0 FreeSans 280 90 0 0 out
port 5 nsew
flabel metal2 s 28557 -656 28613 144 0 FreeSans 280 90 0 0 dout
port 1 nsew
flabel metal2 s 27507 -656 27563 144 0 FreeSans 280 90 0 0 ena
port 3 nsew
flabel metal2 s 30044 -656 30100 144 0 FreeSans 280 90 0 0 stdby
port 4 nsew
flabel metal2 s 89785 42249 89913 43705 0 FreeSans 280 90 0 0 in
port 2 nsew
flabel metal4 s 23284 0 23604 42360 0 FreeSans 2400 90 0 0 vssd1
port 7 nsew
flabel metal4 s 24350 0 24670 42360 0 FreeSans 2400 90 0 0 vssd1
port 7 nsew
flabel metal4 s 31139 0 31459 42360 0 FreeSans 2400 90 0 0 vdda1
port 8 nsew
flabel metal4 s 30310 0 30630 42360 0 FreeSans 2400 90 0 0 vdda1
port 8 nsew
flabel metal4 s 29151 0 29471 42360 0 FreeSans 2400 90 0 0 vccd1
port 9 nsew
flabel metal4 s 27047 0 27367 42360 0 FreeSans 2400 90 0 0 vssa1
port 10 nsew
flabel metal4 s 26142 0 26462 42360 0 FreeSans 2400 90 0 0 vssa1
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 90889 42360
<< end >>
