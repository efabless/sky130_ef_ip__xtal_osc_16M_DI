magic
tech sky130A
magscale 1 2
timestamp 1527871280
<< checkpaint >>
rect 896 -1916 105344 44965
<< metal1 >>
rect 37149 12693 41256 12704
rect 37149 12513 37465 12693
rect 37773 12690 41256 12693
rect 37773 12513 38530 12690
rect 37149 12510 38530 12513
rect 38838 12510 41256 12690
rect 37149 12508 41256 12510
rect 42728 12209 42928 12708
rect 42728 12093 42779 12209
rect 42895 12093 42928 12209
rect 42728 12048 42928 12093
<< via1 >>
rect 41963 23258 42079 23374
rect 43692 23257 43808 23373
rect 37465 12513 37773 12693
rect 38530 12510 38838 12690
rect 41724 12563 41840 12679
rect 44254 12557 44370 12673
rect 42779 12093 42895 12209
<< metal2 >>
rect 2156 27194 2284 43705
rect 103956 27194 104084 43705
rect 2156 26994 42118 27194
rect 41918 23374 42118 26994
rect 41918 23258 41963 23374
rect 42079 23258 42118 23374
rect 41918 23212 42118 23258
rect 43656 26994 104084 27194
rect 43656 23373 43856 26994
rect 43656 23257 43692 23373
rect 43808 23257 43856 23373
rect 43656 23212 43856 23257
rect 37149 12693 39228 12704
rect 37149 12513 37465 12693
rect 37773 12690 39228 12693
rect 37773 12513 38530 12690
rect 37149 12510 38530 12513
rect 38838 12510 39228 12690
rect 37149 12508 39228 12510
rect 41678 12679 41878 12708
rect 41678 12563 41724 12679
rect 41840 12563 41878 12679
rect 44214 12673 44414 12708
rect 41678 0 41878 12563
rect 44214 12557 44254 12673
rect 44370 12557 44414 12673
rect 42728 12209 42928 12330
rect 42728 12093 42779 12209
rect 42895 12093 42928 12209
rect 42728 0 42928 12093
rect 44214 0 44414 12557
rect 41678 -656 41734 0
rect 42728 -656 42784 0
rect 44215 -656 44271 0
<< via2 >>
rect 40319 23324 40375 23380
rect 40399 23324 40455 23380
rect 40479 23324 40535 23380
rect 40559 23324 40615 23380
rect 41224 23324 41280 23380
rect 41304 23324 41360 23380
rect 41384 23324 41440 23380
rect 41464 23324 41520 23380
rect 40319 23235 40375 23291
rect 40399 23235 40455 23291
rect 40479 23235 40535 23291
rect 40559 23235 40615 23291
rect 41224 23230 41280 23286
rect 41304 23230 41360 23286
rect 41384 23230 41440 23286
rect 41464 23230 41520 23286
rect 44487 23324 44543 23380
rect 44567 23324 44623 23380
rect 44647 23324 44703 23380
rect 44727 23324 44783 23380
rect 45316 23324 45372 23380
rect 45396 23324 45452 23380
rect 45476 23324 45532 23380
rect 45556 23324 45612 23380
rect 37469 12620 37525 12676
rect 37549 12620 37605 12676
rect 37629 12620 37685 12676
rect 37709 12620 37765 12676
rect 37469 12531 37525 12587
rect 37549 12531 37605 12587
rect 37629 12531 37685 12587
rect 37709 12531 37765 12587
rect 38534 12620 38590 12676
rect 38614 12620 38670 12676
rect 38694 12620 38750 12676
rect 38774 12620 38830 12676
rect 38534 12526 38590 12582
rect 38614 12526 38670 12582
rect 38694 12526 38750 12582
rect 38774 12526 38830 12582
rect 43340 12598 43396 12654
rect 43420 12598 43476 12654
rect 43500 12598 43556 12654
rect 43580 12598 43636 12654
rect 43340 12509 43396 12565
rect 43420 12509 43476 12565
rect 43500 12509 43556 12565
rect 43580 12509 43636 12565
<< metal3 >>
rect 40225 23384 41850 23412
rect 40225 23320 40315 23384
rect 40379 23320 40395 23384
rect 40459 23320 40475 23384
rect 40539 23320 40555 23384
rect 40619 23320 41220 23384
rect 41284 23320 41300 23384
rect 41364 23320 41380 23384
rect 41444 23320 41460 23384
rect 41524 23320 41850 23384
rect 40225 23295 41850 23320
rect 40225 23231 40315 23295
rect 40379 23231 40395 23295
rect 40459 23231 40475 23295
rect 40539 23231 40555 23295
rect 40619 23290 41850 23295
rect 40619 23231 41220 23290
rect 40225 23226 41220 23231
rect 41284 23226 41300 23290
rect 41364 23226 41380 23290
rect 41444 23226 41460 23290
rect 41524 23226 41850 23290
rect 44227 23384 45855 23412
rect 44227 23320 44483 23384
rect 44547 23320 44563 23384
rect 44627 23320 44643 23384
rect 44707 23320 44723 23384
rect 44787 23320 45312 23384
rect 45376 23320 45392 23384
rect 45456 23320 45472 23384
rect 45536 23320 45552 23384
rect 45616 23320 45855 23384
rect 44227 23287 45855 23320
rect 40225 23210 41850 23226
rect 37375 12680 39000 12708
rect 37375 12616 37465 12680
rect 37529 12616 37545 12680
rect 37609 12616 37625 12680
rect 37689 12616 37705 12680
rect 37769 12616 38530 12680
rect 38594 12616 38610 12680
rect 38674 12616 38690 12680
rect 38754 12616 38770 12680
rect 38834 12616 39000 12680
rect 37375 12591 39000 12616
rect 37375 12527 37465 12591
rect 37529 12527 37545 12591
rect 37609 12527 37625 12591
rect 37689 12527 37705 12591
rect 37769 12586 39000 12591
rect 37769 12527 38530 12586
rect 37375 12522 38530 12527
rect 38594 12522 38610 12586
rect 38674 12522 38690 12586
rect 38754 12522 38770 12586
rect 38834 12522 39000 12586
rect 37375 12506 39000 12522
rect 43246 12658 43830 12686
rect 43246 12594 43336 12658
rect 43400 12594 43416 12658
rect 43480 12594 43496 12658
rect 43560 12594 43576 12658
rect 43640 12594 43830 12658
rect 43246 12569 43830 12594
rect 43246 12505 43336 12569
rect 43400 12505 43416 12569
rect 43480 12505 43496 12569
rect 43560 12505 43576 12569
rect 43640 12505 43830 12569
rect 43246 12484 43830 12505
<< via3 >>
rect 40315 23380 40379 23384
rect 40315 23324 40319 23380
rect 40319 23324 40375 23380
rect 40375 23324 40379 23380
rect 40315 23320 40379 23324
rect 40395 23380 40459 23384
rect 40395 23324 40399 23380
rect 40399 23324 40455 23380
rect 40455 23324 40459 23380
rect 40395 23320 40459 23324
rect 40475 23380 40539 23384
rect 40475 23324 40479 23380
rect 40479 23324 40535 23380
rect 40535 23324 40539 23380
rect 40475 23320 40539 23324
rect 40555 23380 40619 23384
rect 40555 23324 40559 23380
rect 40559 23324 40615 23380
rect 40615 23324 40619 23380
rect 40555 23320 40619 23324
rect 41220 23380 41284 23384
rect 41220 23324 41224 23380
rect 41224 23324 41280 23380
rect 41280 23324 41284 23380
rect 41220 23320 41284 23324
rect 41300 23380 41364 23384
rect 41300 23324 41304 23380
rect 41304 23324 41360 23380
rect 41360 23324 41364 23380
rect 41300 23320 41364 23324
rect 41380 23380 41444 23384
rect 41380 23324 41384 23380
rect 41384 23324 41440 23380
rect 41440 23324 41444 23380
rect 41380 23320 41444 23324
rect 41460 23380 41524 23384
rect 41460 23324 41464 23380
rect 41464 23324 41520 23380
rect 41520 23324 41524 23380
rect 41460 23320 41524 23324
rect 40315 23291 40379 23295
rect 40315 23235 40319 23291
rect 40319 23235 40375 23291
rect 40375 23235 40379 23291
rect 40315 23231 40379 23235
rect 40395 23291 40459 23295
rect 40395 23235 40399 23291
rect 40399 23235 40455 23291
rect 40455 23235 40459 23291
rect 40395 23231 40459 23235
rect 40475 23291 40539 23295
rect 40475 23235 40479 23291
rect 40479 23235 40535 23291
rect 40535 23235 40539 23291
rect 40475 23231 40539 23235
rect 40555 23291 40619 23295
rect 40555 23235 40559 23291
rect 40559 23235 40615 23291
rect 40615 23235 40619 23291
rect 40555 23231 40619 23235
rect 41220 23286 41284 23290
rect 41220 23230 41224 23286
rect 41224 23230 41280 23286
rect 41280 23230 41284 23286
rect 41220 23226 41284 23230
rect 41300 23286 41364 23290
rect 41300 23230 41304 23286
rect 41304 23230 41360 23286
rect 41360 23230 41364 23286
rect 41300 23226 41364 23230
rect 41380 23286 41444 23290
rect 41380 23230 41384 23286
rect 41384 23230 41440 23286
rect 41440 23230 41444 23286
rect 41380 23226 41444 23230
rect 41460 23286 41524 23290
rect 41460 23230 41464 23286
rect 41464 23230 41520 23286
rect 41520 23230 41524 23286
rect 41460 23226 41524 23230
rect 44483 23380 44547 23384
rect 44483 23324 44487 23380
rect 44487 23324 44543 23380
rect 44543 23324 44547 23380
rect 44483 23320 44547 23324
rect 44563 23380 44627 23384
rect 44563 23324 44567 23380
rect 44567 23324 44623 23380
rect 44623 23324 44627 23380
rect 44563 23320 44627 23324
rect 44643 23380 44707 23384
rect 44643 23324 44647 23380
rect 44647 23324 44703 23380
rect 44703 23324 44707 23380
rect 44643 23320 44707 23324
rect 44723 23380 44787 23384
rect 44723 23324 44727 23380
rect 44727 23324 44783 23380
rect 44783 23324 44787 23380
rect 44723 23320 44787 23324
rect 45312 23380 45376 23384
rect 45312 23324 45316 23380
rect 45316 23324 45372 23380
rect 45372 23324 45376 23380
rect 45312 23320 45376 23324
rect 45392 23380 45456 23384
rect 45392 23324 45396 23380
rect 45396 23324 45452 23380
rect 45452 23324 45456 23380
rect 45392 23320 45456 23324
rect 45472 23380 45536 23384
rect 45472 23324 45476 23380
rect 45476 23324 45532 23380
rect 45532 23324 45536 23380
rect 45472 23320 45536 23324
rect 45552 23380 45616 23384
rect 45552 23324 45556 23380
rect 45556 23324 45612 23380
rect 45612 23324 45616 23380
rect 45552 23320 45616 23324
rect 37465 12676 37529 12680
rect 37465 12620 37469 12676
rect 37469 12620 37525 12676
rect 37525 12620 37529 12676
rect 37465 12616 37529 12620
rect 37545 12676 37609 12680
rect 37545 12620 37549 12676
rect 37549 12620 37605 12676
rect 37605 12620 37609 12676
rect 37545 12616 37609 12620
rect 37625 12676 37689 12680
rect 37625 12620 37629 12676
rect 37629 12620 37685 12676
rect 37685 12620 37689 12676
rect 37625 12616 37689 12620
rect 37705 12676 37769 12680
rect 37705 12620 37709 12676
rect 37709 12620 37765 12676
rect 37765 12620 37769 12676
rect 37705 12616 37769 12620
rect 38530 12676 38594 12680
rect 38530 12620 38534 12676
rect 38534 12620 38590 12676
rect 38590 12620 38594 12676
rect 38530 12616 38594 12620
rect 38610 12676 38674 12680
rect 38610 12620 38614 12676
rect 38614 12620 38670 12676
rect 38670 12620 38674 12676
rect 38610 12616 38674 12620
rect 38690 12676 38754 12680
rect 38690 12620 38694 12676
rect 38694 12620 38750 12676
rect 38750 12620 38754 12676
rect 38690 12616 38754 12620
rect 38770 12676 38834 12680
rect 38770 12620 38774 12676
rect 38774 12620 38830 12676
rect 38830 12620 38834 12676
rect 38770 12616 38834 12620
rect 37465 12587 37529 12591
rect 37465 12531 37469 12587
rect 37469 12531 37525 12587
rect 37525 12531 37529 12587
rect 37465 12527 37529 12531
rect 37545 12587 37609 12591
rect 37545 12531 37549 12587
rect 37549 12531 37605 12587
rect 37605 12531 37609 12587
rect 37545 12527 37609 12531
rect 37625 12587 37689 12591
rect 37625 12531 37629 12587
rect 37629 12531 37685 12587
rect 37685 12531 37689 12587
rect 37625 12527 37689 12531
rect 37705 12587 37769 12591
rect 37705 12531 37709 12587
rect 37709 12531 37765 12587
rect 37765 12531 37769 12587
rect 37705 12527 37769 12531
rect 38530 12582 38594 12586
rect 38530 12526 38534 12582
rect 38534 12526 38590 12582
rect 38590 12526 38594 12582
rect 38530 12522 38594 12526
rect 38610 12582 38674 12586
rect 38610 12526 38614 12582
rect 38614 12526 38670 12582
rect 38670 12526 38674 12582
rect 38610 12522 38674 12526
rect 38690 12582 38754 12586
rect 38690 12526 38694 12582
rect 38694 12526 38750 12582
rect 38750 12526 38754 12582
rect 38690 12522 38754 12526
rect 38770 12582 38834 12586
rect 38770 12526 38774 12582
rect 38774 12526 38830 12582
rect 38830 12526 38834 12582
rect 38770 12522 38834 12526
rect 43336 12654 43400 12658
rect 43336 12598 43340 12654
rect 43340 12598 43396 12654
rect 43396 12598 43400 12654
rect 43336 12594 43400 12598
rect 43416 12654 43480 12658
rect 43416 12598 43420 12654
rect 43420 12598 43476 12654
rect 43476 12598 43480 12654
rect 43416 12594 43480 12598
rect 43496 12654 43560 12658
rect 43496 12598 43500 12654
rect 43500 12598 43556 12654
rect 43556 12598 43560 12654
rect 43496 12594 43560 12598
rect 43576 12654 43640 12658
rect 43576 12598 43580 12654
rect 43580 12598 43636 12654
rect 43636 12598 43640 12654
rect 43576 12594 43640 12598
rect 43336 12565 43400 12569
rect 43336 12509 43340 12565
rect 43340 12509 43396 12565
rect 43396 12509 43400 12565
rect 43336 12505 43400 12509
rect 43416 12565 43480 12569
rect 43416 12509 43420 12565
rect 43420 12509 43476 12565
rect 43476 12509 43480 12565
rect 43416 12505 43480 12509
rect 43496 12565 43560 12569
rect 43496 12509 43500 12565
rect 43500 12509 43556 12565
rect 43556 12509 43560 12565
rect 43496 12505 43560 12509
rect 43576 12565 43640 12569
rect 43576 12509 43580 12565
rect 43580 12509 43636 12565
rect 43636 12509 43640 12565
rect 43576 12505 43640 12509
<< metal4 >>
rect 37455 12680 37775 42360
rect 37455 12616 37465 12680
rect 37529 12616 37545 12680
rect 37609 12616 37625 12680
rect 37689 12616 37705 12680
rect 37769 12616 37775 12680
rect 37455 12591 37775 12616
rect 37455 12527 37465 12591
rect 37529 12527 37545 12591
rect 37609 12527 37625 12591
rect 37689 12527 37705 12591
rect 37769 12527 37775 12591
rect 37455 0 37775 12527
rect 38521 12680 38841 42360
rect 38521 12616 38530 12680
rect 38594 12616 38610 12680
rect 38674 12616 38690 12680
rect 38754 12616 38770 12680
rect 38834 12616 38841 12680
rect 38521 12586 38841 12616
rect 38521 12522 38530 12586
rect 38594 12522 38610 12586
rect 38674 12522 38690 12586
rect 38754 12522 38770 12586
rect 38834 12522 38841 12586
rect 38521 0 38841 12522
rect 40313 23384 40633 42360
rect 40313 23320 40315 23384
rect 40379 23320 40395 23384
rect 40459 23320 40475 23384
rect 40539 23320 40555 23384
rect 40619 23320 40633 23384
rect 40313 23295 40633 23320
rect 40313 23231 40315 23295
rect 40379 23231 40395 23295
rect 40459 23231 40475 23295
rect 40539 23231 40555 23295
rect 40619 23231 40633 23295
rect 40313 0 40633 23231
rect 41218 23384 41538 42360
rect 41218 23320 41220 23384
rect 41284 23320 41300 23384
rect 41364 23320 41380 23384
rect 41444 23320 41460 23384
rect 41524 23320 41538 23384
rect 41218 23290 41538 23320
rect 41218 23226 41220 23290
rect 41284 23226 41300 23290
rect 41364 23226 41380 23290
rect 41444 23226 41460 23290
rect 41524 23226 41538 23290
rect 41218 0 41538 23226
rect 43322 12658 43642 42360
rect 43322 12594 43336 12658
rect 43400 12594 43416 12658
rect 43480 12594 43496 12658
rect 43560 12594 43576 12658
rect 43640 12594 43642 12658
rect 43322 12569 43642 12594
rect 43322 12505 43336 12569
rect 43400 12505 43416 12569
rect 43480 12505 43496 12569
rect 43560 12505 43576 12569
rect 43640 12505 43642 12569
rect 43322 0 43642 12505
rect 44481 23384 44801 42360
rect 44481 23320 44483 23384
rect 44547 23320 44563 23384
rect 44627 23320 44643 23384
rect 44707 23320 44723 23384
rect 44787 23320 44801 23384
rect 44481 0 44801 23320
rect 45310 23384 45630 42360
rect 45310 23320 45312 23384
rect 45376 23320 45392 23384
rect 45456 23320 45472 23384
rect 45536 23320 45552 23384
rect 45616 23320 45630 23384
rect 45310 0 45630 23320
use sky130_ef_ip__xtal_osc_16M  sky130_ef_ip__xtal_osc_16M_0
timestamp 1527871280
transform 0 1 42640 -1 0 25872
box 2460 -2440 13388 3256
<< labels >>
flabel metal2 s 42728 -656 42784 144 0 FreeSans 280 90 0 0 dout
port 1 nsew
flabel metal2 s 41678 -656 41734 144 0 FreeSans 280 90 0 0 ena
port 4 nsew
flabel metal2 s 44215 -656 44271 144 0 FreeSans 280 90 0 0 stdby
port 5 nsew
flabel metal2 s 2156 42249 2284 43705 0 FreeSans 280 90 0 0 out
port 3 nsew
flabel metal2 s 103956 42249 104084 43705 0 FreeSans 280 90 0 0 in
port 2 nsew
flabel metal4 s 37455 0 37775 42360 0 FreeSans 2400 90 0 0 vssd1
port 7 nsew
flabel metal4 s 38521 0 38841 42360 0 FreeSans 2400 90 0 0 vssd1
port 7 nsew
flabel metal4 s 45310 0 45630 42360 0 FreeSans 2400 90 0 0 vdda1
port 8 nsew
flabel metal4 s 44481 0 44801 42360 0 FreeSans 2400 90 0 0 vdda1
port 8 nsew
flabel metal4 s 43322 0 43642 42360 0 FreeSans 2400 90 0 0 vccd1
port 9 nsew
flabel metal4 s 41218 0 41538 42360 0 FreeSans 2400 90 0 0 vssa1
port 10 nsew
flabel metal4 s 40313 0 40633 42360 0 FreeSans 2400 90 0 0 vssa1
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 105060 42360
<< end >>
